* Tue Aug 10 11:21:07 CEST 2004
.subckt nd4_x1 a b c d vdd vss z 
*SPICE circuit <nd4_x1> from XCircuit v3.10

m1 n1 a vss vss n w=32u l=2.3636u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m2 n2 b n1 vss n w=32u l=2.3636u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m3 n3 c n2 vss n w=32u l=2.3636u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m4 z d n3 vss n w=32u l=2.3636u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m5 z a vdd vdd p w=27u l=2.3636u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
m6 z b vdd vdd p w=27u l=2.3636u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
m7 z c vdd vdd p w=27u l=2.3636u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
m8 z d vdd vdd p w=27u l=2.3636u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
.ends
