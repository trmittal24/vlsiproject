* Thu Jan 11 12:51:16 CET 2007
.subckt mxi2v2x1 a0 a1 s vdd vss z
*SPICE circuit <mxi2v2x1> from XCircuit v3.20

m1 a0n a0 vdd vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m2 a1n a1 vdd vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m3 z sn a1n vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m4 a0n s z vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m5 sn s vdd vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m6 a1n a1 vss vss n w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m7 z sn a0n vss n w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m8 a1n s z vss n w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m9 a0n a0 vss vss n w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m10 sn s vss vss n w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
.ends
