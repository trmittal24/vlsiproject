* Spice description of vfeed1
* Spice driver version 134999461
* Date 22/07/2007 at 11:00:16
* vsxlib 0.13um values
.subckt vfeed1 vdd vss
.ends
