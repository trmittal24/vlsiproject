* Sat Apr  9 11:31:05 CEST 2005
.subckt nr3v0x4 a b c vdd vss z 
*SPICE circuit <nr3v0x4> from XCircuit v3.20

m1 z a vss vss n w=24u l=2u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m2 z c vss vss n w=24u l=2u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m3 n1 a vdd vdd p w=132u l=2u ad='132u*5u+12p' as='132u*5u+12p' pd='132u*2+14u' ps='132u*2+14u'
m4 n2 b n1 vdd p w=132u l=2u ad='132u*5u+12p' as='132u*5u+12p' pd='132u*2+14u' ps='132u*2+14u'
m5 z b vss vss n w=24u l=2u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m6 z c n2 vdd p w=132u l=2u ad='132u*5u+12p' as='132u*5u+12p' pd='132u*2+14u' ps='132u*2+14u'
.ends
