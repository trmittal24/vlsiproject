* Fri Dec  8 16:10:46 CET 2006
.subckt cgi2bv0x05 a b c vdd vss z
*SPICE circuit <cgi2bv0x05> from XCircuit v3.20

m1 bn b vdd vdd p w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m2 bn b vss vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m3 n1 bn vdd vdd p w=16u l=2.3636u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m4 n1 a vdd vdd p w=16u l=2.3636u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m5 z c n1 vdd p w=16u l=2.3636u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m6 n2 a vdd vdd p w=16u l=2.3636u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m7 z bn n2 vdd p w=16u l=2.3636u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m8 n3 bn vss vss n w=7u l=2.3636u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m9 n3 a vss vss n w=7u l=2.3636u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m10 n4 a vss vss n w=7u l=2.3636u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m11 z bn n4 vss n w=7u l=2.3636u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m12 z c n3 vss n w=7u l=2.3636u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
.ends
