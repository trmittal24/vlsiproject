* Spice description of o2_x2
* Spice driver version 134999461
* Date 31/05/2007 at 10:39:28
* ssxlib 0.13um values
.subckt o2_x2 i0 i1 q vdd vss
Mtr_00001 q     sig1  vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00002 sig1  i0    vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00003 vss   i1    sig1  vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00004 sig6  i1    sig1  vdd p  L=0.12U  W=1.595U AS=0.422675P AD=0.422675P PS=3.72U   PD=3.72U
Mtr_00005 vdd   i0    sig6  vdd p  L=0.12U  W=1.595U AS=0.422675P AD=0.422675P PS=3.72U   PD=3.72U
Mtr_00006 q     sig1  vdd   vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
C3  i0    vss   0.927f
C4  i1    vss   0.646f
C5  q     vss   0.900f
C1  sig1  vss   0.748f
.ends
