* Spice description of vfeed4
* Spice driver version 134999461
* Date 31/05/2007 at 21:36:02
* vxlib 0.13um values
.subckt vfeed4 vdd vss
.ends
