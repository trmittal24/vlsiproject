magic
tech scmos
timestamp 1523104733
<< polysilicon >>
rect 815 304 817 313
rect 1024 148 1026 156
rect 1041 147 1043 156
rect 1048 149 1050 162
<< metal1 >>
rect 841 506 885 510
rect 839 421 875 425
rect 119 362 157 366
rect 152 245 157 362
rect 839 343 854 347
rect 858 343 859 347
rect 1050 310 1051 314
rect 813 294 817 300
rect 1041 295 1042 299
rect 1024 271 1025 275
rect 697 247 857 250
rect 152 241 425 245
rect 675 228 720 230
rect 675 222 721 228
rect 676 220 721 222
rect 430 195 630 198
rect 676 162 727 164
rect 676 155 866 162
rect 1022 160 1025 271
rect 1039 160 1042 295
rect 1048 166 1051 310
rect 1050 162 1051 166
rect 680 149 866 155
rect 817 144 830 149
rect 972 144 985 152
rect 461 98 464 129
rect 810 102 952 106
rect 818 80 831 88
rect 969 80 982 88
<< metal2 >>
rect 889 506 890 510
rect 879 421 880 425
rect 654 367 665 370
rect 381 362 402 366
rect 641 362 665 367
rect 33 195 106 198
rect 399 199 402 362
rect 654 360 665 362
rect 833 343 841 347
rect 858 343 859 346
rect 814 294 817 295
rect 328 195 402 199
rect 693 243 697 246
rect 814 243 817 290
rect 856 275 859 343
rect 877 299 880 421
rect 887 314 890 506
rect 887 310 1046 314
rect 877 295 1037 299
rect 856 271 1020 275
rect 425 199 429 241
rect 461 240 697 243
rect 753 240 817 243
rect 461 133 464 240
rect 753 203 756 240
rect 858 202 861 247
rect 754 191 810 194
rect 807 123 810 191
rect 952 109 981 113
rect 952 107 957 109
<< metal3 >>
rect 653 359 666 371
rect 108 263 119 264
rect 654 263 666 359
rect 107 253 666 263
rect 108 204 119 253
rect 104 202 122 204
rect 104 190 106 202
rect 120 190 122 202
rect 104 188 122 190
<< polycontact >>
rect 813 300 817 304
rect 1046 162 1050 166
rect 1022 156 1026 160
rect 1039 156 1043 160
<< m2contact >>
rect 885 506 889 510
rect 875 421 879 425
rect 854 343 858 347
rect 1046 310 1050 314
rect 1037 295 1041 299
rect 813 290 817 294
rect 1020 271 1024 275
rect 693 246 697 250
rect 857 247 861 251
rect 425 241 430 246
rect 753 199 757 203
rect 425 195 430 199
rect 858 198 862 202
rect 750 191 754 195
rect 461 129 465 133
rect 807 119 811 123
rect 981 109 985 113
rect 952 102 957 107
rect 461 94 465 98
<< m3contact >>
rect 106 190 120 202
<< psubstratepcontact >>
rect 654 360 665 370
use totdiff3  totdiff3_0
timestamp 1523087024
transform 1 0 -569 0 1 937
box 507 -672 1412 -374
use dfnt1v0x2  dfnt1v0x2_1
timestamp 1523100110
transform -1 0 864 0 -1 232
box -4 -4 148 76
use ../../../../prac/counter  counter_0
timestamp 1523087024
transform 1 0 608 0 1 76
box -608 -76 216 157
use or3v0x3  or3v0x3_0
timestamp 1523091398
transform 1 0 979 0 1 80
box -4 -4 84 76
<< end >>
