* Mon Aug 16 14:10:58 CEST 2004
.subckt iv1v0x4 a vdd vss z 
*SPICE circuit <iv1v0x4> from XCircuit v3.10

m1 z a vss vss n w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m2 z a vdd vdd p w=56u l=2.3636u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
.ends
