* Thu Sep  1 18:58:48 CEST 2005
.subckt nr2v1x4 a b vdd vss z 
*SPICE circuit <nr2v1x4> from XCircuit v3.20

m1 z a vss vss n w=53u l=2.3636u ad='53u*5u+12p' as='53u*5u+12p' pd='53u*2+14u' ps='53u*2+14u'
m2 n1 a vdd vdd p w=108u l=2.3636u ad='108u*5u+12p' as='108u*5u+12p' pd='108u*2+14u' ps='108u*2+14u'
m3 z b vss vss n w=53u l=2.3636u ad='53u*5u+12p' as='53u*5u+12p' pd='53u*2+14u' ps='53u*2+14u'
m4 z b n1 vdd p w=108u l=2.3636u ad='108u*5u+12p' as='108u*5u+12p' pd='108u*2+14u' ps='108u*2+14u'
.ends
