magic
tech scmos
timestamp 1522862826
<< pwell >>
rect -139 0 152 36
<< nwell >>
rect -139 36 152 80
<< polysilicon >>
rect -115 70 -113 74
rect -105 70 -103 74
rect -90 70 -88 74
rect -80 70 -78 74
rect -50 70 -48 74
rect -40 70 -38 74
rect -30 70 -28 74
rect -20 70 -18 74
rect -10 70 -8 74
rect 13 70 15 74
rect -64 63 -58 64
rect -70 55 -68 60
rect -64 59 -63 63
rect -59 59 -58 63
rect -64 58 -58 59
rect -60 55 -58 58
rect 59 72 115 74
rect 59 64 61 72
rect 69 64 71 68
rect 79 64 81 68
rect 86 64 88 72
rect 96 64 98 68
rect 103 64 105 68
rect 23 56 25 61
rect 42 58 44 63
rect 49 58 51 63
rect -115 39 -113 42
rect -105 39 -103 42
rect -90 39 -88 42
rect -80 39 -78 42
rect -126 38 -84 39
rect -126 34 -125 38
rect -121 37 -84 38
rect -121 34 -114 37
rect -126 33 -114 34
rect -126 30 -124 33
rect -116 30 -114 33
rect -96 30 -94 37
rect -86 30 -84 37
rect -80 38 -74 39
rect -80 34 -79 38
rect -75 34 -74 38
rect -70 37 -68 42
rect -60 37 -58 42
rect -50 39 -48 42
rect -40 39 -38 42
rect -30 39 -28 42
rect -50 38 -38 39
rect -70 35 -55 37
rect -80 33 -74 34
rect -76 30 -74 33
rect -69 30 -67 35
rect -57 30 -55 35
rect -50 34 -49 38
rect -45 37 -38 38
rect -34 38 -28 39
rect -45 34 -44 37
rect -50 33 -44 34
rect -34 34 -33 38
rect -29 34 -28 38
rect -34 33 -28 34
rect -20 39 -18 42
rect -10 39 -8 42
rect -20 38 -8 39
rect -20 34 -13 38
rect -9 34 -8 38
rect -20 33 -8 34
rect -50 30 -48 33
rect -20 30 -18 33
rect -10 30 -8 33
rect 13 38 15 42
rect 23 39 25 42
rect 23 38 38 39
rect 13 37 19 38
rect 23 37 33 38
rect 13 33 14 37
rect 18 33 19 37
rect 13 32 19 33
rect 31 34 33 37
rect 37 34 38 38
rect 31 33 38 34
rect -126 15 -124 19
rect -116 8 -114 13
rect -96 11 -94 16
rect -86 11 -84 16
rect -76 6 -74 11
rect -69 6 -67 11
rect 13 28 15 32
rect 31 30 33 33
rect -20 12 -18 16
rect -10 12 -8 16
rect 42 23 44 52
rect 49 48 51 52
rect 49 47 55 48
rect 49 43 50 47
rect 54 43 55 47
rect 49 42 55 43
rect 59 38 61 52
rect 49 36 61 38
rect 49 23 51 36
rect 69 33 71 52
rect 79 48 81 58
rect 75 47 81 48
rect 75 43 76 47
rect 80 43 81 47
rect 75 42 81 43
rect 69 32 75 33
rect 55 31 61 32
rect 55 27 56 31
rect 60 27 61 31
rect 55 26 61 27
rect 59 23 61 26
rect 69 28 70 32
rect 74 28 75 32
rect 69 27 75 28
rect 69 23 71 27
rect 79 23 81 42
rect 86 38 88 58
rect 113 62 115 72
rect 133 63 135 68
rect 96 48 98 51
rect 92 47 98 48
rect 92 43 93 47
rect 97 43 98 47
rect 92 42 98 43
rect 103 39 105 51
rect 113 48 115 51
rect 133 49 135 53
rect 126 48 135 49
rect 113 46 121 48
rect 119 39 121 46
rect 126 44 127 48
rect 131 44 135 48
rect 126 43 135 44
rect 103 38 109 39
rect 86 36 98 38
rect 86 31 92 32
rect 86 27 87 31
rect 91 27 92 31
rect 86 26 92 27
rect 86 23 88 26
rect 96 23 98 36
rect 103 34 104 38
rect 108 34 109 38
rect 103 33 109 34
rect 119 38 125 39
rect 119 34 120 38
rect 124 34 125 38
rect 119 33 125 34
rect 103 23 105 33
rect 123 30 125 33
rect 133 30 135 43
rect 31 18 33 23
rect 123 19 125 24
rect 133 18 135 23
rect -57 6 -55 11
rect -50 6 -48 11
rect 13 11 15 14
rect 42 11 44 17
rect 49 12 51 17
rect 13 9 44 11
rect 59 8 61 17
rect 69 12 71 17
rect 79 12 81 17
rect 86 8 88 17
rect 96 12 98 17
rect 103 12 105 17
rect 59 6 88 8
<< ndiffusion >>
rect -133 24 -126 30
rect -133 20 -132 24
rect -128 20 -126 24
rect -133 19 -126 20
rect -124 29 -116 30
rect -124 25 -122 29
rect -118 25 -116 29
rect -124 19 -116 25
rect -121 13 -116 19
rect -114 18 -107 30
rect -114 14 -112 18
rect -108 14 -107 18
rect -103 29 -96 30
rect -103 25 -102 29
rect -98 25 -96 29
rect -103 22 -96 25
rect -103 18 -102 22
rect -98 18 -96 22
rect -103 16 -96 18
rect -94 29 -86 30
rect -94 25 -92 29
rect -88 25 -86 29
rect -94 16 -86 25
rect -84 29 -76 30
rect -84 25 -82 29
rect -78 25 -76 29
rect -84 22 -76 25
rect -84 18 -82 22
rect -78 18 -76 22
rect -84 16 -76 18
rect -114 13 -107 14
rect -81 11 -76 16
rect -74 11 -69 30
rect -67 12 -57 30
rect -67 11 -64 12
rect -65 8 -64 11
rect -60 11 -57 12
rect -55 11 -50 30
rect -48 23 -43 30
rect -48 22 -41 23
rect -48 18 -46 22
rect -42 18 -41 22
rect -48 17 -41 18
rect -48 11 -43 17
rect -27 21 -20 30
rect -27 17 -26 21
rect -22 17 -20 21
rect -27 16 -20 17
rect -18 29 -10 30
rect -18 25 -16 29
rect -12 25 -10 29
rect -18 22 -10 25
rect -18 18 -16 22
rect -12 18 -10 22
rect -18 16 -10 18
rect -8 21 -1 30
rect 24 29 31 30
rect 6 27 13 28
rect 6 23 7 27
rect 11 23 13 27
rect 6 22 13 23
rect -8 17 -6 21
rect -2 17 -1 21
rect -8 16 -1 17
rect 8 14 13 22
rect 15 20 20 28
rect 24 25 25 29
rect 29 25 31 29
rect 24 24 31 25
rect 26 23 31 24
rect 33 23 40 30
rect 116 29 123 30
rect 116 25 117 29
rect 121 25 123 29
rect 116 24 123 25
rect 125 29 133 30
rect 125 25 127 29
rect 131 25 133 29
rect 125 24 133 25
rect 15 19 22 20
rect 15 15 17 19
rect 21 15 22 19
rect 35 22 42 23
rect 35 18 36 22
rect 40 18 42 22
rect 35 17 42 18
rect 44 17 49 23
rect 51 22 59 23
rect 51 18 53 22
rect 57 18 59 22
rect 51 17 59 18
rect 61 22 69 23
rect 61 18 63 22
rect 67 18 69 22
rect 61 17 69 18
rect 71 22 79 23
rect 71 18 73 22
rect 77 18 79 22
rect 71 17 79 18
rect 81 17 86 23
rect 88 22 96 23
rect 88 18 90 22
rect 94 18 96 22
rect 88 17 96 18
rect 98 17 103 23
rect 105 22 112 23
rect 105 18 107 22
rect 111 18 112 22
rect 127 23 133 24
rect 135 29 142 30
rect 135 25 137 29
rect 141 25 142 29
rect 135 23 142 25
rect 105 17 112 18
rect 15 14 22 15
rect -60 8 -59 11
rect -65 7 -59 8
<< pdiffusion >>
rect -122 69 -115 70
rect -122 65 -121 69
rect -117 65 -115 69
rect -122 62 -115 65
rect -122 58 -121 62
rect -117 58 -115 62
rect -122 42 -115 58
rect -113 54 -105 70
rect -113 50 -111 54
rect -107 50 -105 54
rect -113 47 -105 50
rect -113 43 -111 47
rect -107 43 -105 47
rect -113 42 -105 43
rect -103 69 -90 70
rect -103 65 -99 69
rect -95 65 -90 69
rect -103 62 -90 65
rect -103 58 -99 62
rect -95 58 -90 62
rect -103 42 -90 58
rect -88 62 -80 70
rect -88 58 -86 62
rect -82 58 -80 62
rect -88 55 -80 58
rect -88 51 -86 55
rect -82 51 -80 55
rect -88 42 -80 51
rect -78 55 -73 70
rect -55 55 -50 70
rect -78 54 -70 55
rect -78 50 -76 54
rect -72 50 -70 54
rect -78 47 -70 50
rect -78 43 -76 47
rect -72 43 -70 47
rect -78 42 -70 43
rect -68 47 -60 55
rect -68 43 -66 47
rect -62 43 -60 47
rect -68 42 -60 43
rect -58 54 -50 55
rect -58 50 -56 54
rect -52 50 -50 54
rect -58 42 -50 50
rect -48 63 -40 70
rect -48 59 -46 63
rect -42 59 -40 63
rect -48 47 -40 59
rect -48 43 -46 47
rect -42 43 -40 47
rect -48 42 -40 43
rect -38 62 -30 70
rect -38 58 -36 62
rect -32 58 -30 62
rect -38 55 -30 58
rect -38 51 -36 55
rect -32 51 -30 55
rect -38 42 -30 51
rect -28 54 -20 70
rect -28 50 -26 54
rect -22 50 -20 54
rect -28 47 -20 50
rect -28 43 -26 47
rect -22 43 -20 47
rect -28 42 -20 43
rect -18 69 -10 70
rect -18 65 -16 69
rect -12 65 -10 69
rect -18 62 -10 65
rect -18 58 -16 62
rect -12 58 -10 62
rect -18 42 -10 58
rect -8 55 -3 70
rect 8 56 13 70
rect -8 54 -1 55
rect -8 50 -6 54
rect -2 50 -1 54
rect -8 47 -1 50
rect -8 43 -6 47
rect -2 43 -1 47
rect -8 42 -1 43
rect 6 54 13 56
rect 6 50 7 54
rect 11 50 13 54
rect 6 47 13 50
rect 6 43 7 47
rect 11 43 13 47
rect 6 42 13 43
rect 15 69 22 70
rect 15 65 17 69
rect 21 65 22 69
rect 15 64 22 65
rect 15 56 21 64
rect 54 58 59 64
rect 34 57 42 58
rect 15 55 23 56
rect 15 51 17 55
rect 21 51 23 55
rect 15 42 23 51
rect 25 48 30 56
rect 34 53 35 57
rect 39 53 42 57
rect 34 52 42 53
rect 44 52 49 58
rect 51 57 59 58
rect 51 53 53 57
rect 57 53 59 57
rect 51 52 59 53
rect 61 57 69 64
rect 61 53 63 57
rect 67 53 69 57
rect 61 52 69 53
rect 71 63 79 64
rect 71 59 73 63
rect 77 59 79 63
rect 71 58 79 59
rect 81 58 86 64
rect 88 63 96 64
rect 88 59 90 63
rect 94 59 96 63
rect 88 58 96 59
rect 71 52 77 58
rect 25 47 32 48
rect 25 43 27 47
rect 31 43 32 47
rect 25 42 32 43
rect 91 51 96 58
rect 98 51 103 64
rect 105 62 110 64
rect 126 62 133 63
rect 105 61 113 62
rect 105 57 107 61
rect 111 57 113 61
rect 105 51 113 57
rect 115 57 120 62
rect 126 58 127 62
rect 131 58 133 62
rect 115 56 122 57
rect 115 52 117 56
rect 121 52 122 56
rect 126 53 133 58
rect 135 59 140 63
rect 135 58 142 59
rect 135 54 137 58
rect 141 54 142 58
rect 135 53 142 54
rect 115 51 122 52
<< metal1 >>
rect -137 72 150 76
rect -137 68 -131 72
rect -127 69 -66 72
rect -127 68 -121 69
rect -117 68 -99 69
rect -121 62 -117 65
rect -100 65 -99 68
rect -95 68 -66 69
rect -62 69 31 72
rect -62 68 -16 69
rect -95 65 -94 68
rect -100 62 -94 65
rect -12 68 17 69
rect -100 58 -99 62
rect -95 58 -94 62
rect -86 62 -63 63
rect -82 59 -63 62
rect -59 59 -46 63
rect -42 59 -41 63
rect -37 62 -32 63
rect -121 57 -117 58
rect -86 55 -82 58
rect -112 50 -111 54
rect -107 51 -86 54
rect -37 58 -36 62
rect -37 55 -32 58
rect -16 62 -12 65
rect -16 57 -12 58
rect 21 68 31 69
rect 35 68 41 72
rect 45 68 122 72
rect 126 68 150 72
rect 17 55 21 65
rect -37 54 -36 55
rect -107 50 -82 51
rect -77 50 -76 54
rect -72 50 -56 54
rect -52 51 -36 54
rect -52 50 -32 51
rect -27 54 -22 55
rect -27 50 -26 54
rect -112 47 -107 50
rect -133 39 -129 47
rect -112 43 -111 47
rect -77 47 -72 50
rect -27 47 -22 50
rect -6 54 -1 55
rect -2 50 -1 54
rect -6 47 -1 50
rect -77 46 -76 47
rect -112 42 -107 43
rect -101 43 -76 46
rect -101 42 -72 43
rect -67 43 -66 47
rect -62 43 -61 47
rect -133 38 -121 39
rect -133 34 -125 38
rect -133 33 -121 34
rect -112 29 -108 42
rect -101 29 -97 42
rect -67 38 -61 43
rect -47 43 -46 47
rect -42 46 -41 47
rect -42 43 -32 46
rect -27 43 -26 47
rect -22 43 -6 47
rect -2 43 -1 47
rect 6 54 11 55
rect 6 50 7 54
rect 35 57 39 68
rect 73 63 77 68
rect 73 58 77 59
rect 85 59 90 63
rect 94 59 95 63
rect 106 61 112 68
rect 63 57 67 58
rect 35 52 39 53
rect 42 53 53 57
rect 57 53 58 57
rect 17 50 21 51
rect 6 47 11 50
rect 6 43 7 47
rect 11 43 19 46
rect -47 42 -32 43
rect -36 38 -32 42
rect -123 25 -122 29
rect -118 25 -108 29
rect -103 25 -102 29
rect -98 25 -97 29
rect -93 34 -79 38
rect -75 34 -49 38
rect -45 34 -42 38
rect -36 34 -33 38
rect -29 34 -28 38
rect -93 29 -87 34
rect -46 30 -42 34
rect -23 30 -19 43
rect 6 42 19 43
rect 25 43 27 47
rect 31 43 32 47
rect -14 38 -1 39
rect -14 34 -13 38
rect -9 34 -1 38
rect 6 34 10 42
rect 25 37 29 43
rect 42 38 46 53
rect 63 47 67 53
rect 49 43 50 47
rect -5 31 10 34
rect 13 33 14 37
rect 18 33 29 37
rect 32 34 33 38
rect 37 34 48 38
rect -93 25 -92 29
rect -88 25 -87 29
rect -82 29 -78 30
rect -46 29 -12 30
rect -46 26 -16 29
rect -132 24 -128 25
rect -132 12 -128 20
rect -103 22 -97 25
rect -82 22 -78 25
rect -5 25 -1 31
rect 6 28 10 31
rect 25 29 29 33
rect 6 27 11 28
rect -16 22 -12 25
rect 6 23 7 27
rect 25 24 29 25
rect 6 22 11 23
rect 36 22 40 23
rect -112 18 -108 19
rect -103 18 -102 22
rect -98 18 -82 22
rect -78 18 -46 22
rect -42 18 -40 22
rect -26 21 -22 22
rect -112 12 -108 14
rect -16 17 -12 18
rect -7 17 -6 21
rect -2 17 -1 21
rect -26 12 -22 17
rect -7 12 -1 17
rect 17 19 21 20
rect 17 12 21 15
rect 44 22 48 34
rect 54 32 58 47
rect 63 43 76 47
rect 80 43 81 47
rect 54 31 60 32
rect 54 27 56 31
rect 54 26 60 27
rect 63 22 67 43
rect 85 40 89 59
rect 106 57 107 61
rect 111 57 112 61
rect 126 62 132 68
rect 126 58 127 62
rect 131 58 132 62
rect 137 58 141 59
rect 117 56 121 57
rect 80 36 89 40
rect 93 52 117 54
rect 93 50 121 52
rect 93 47 97 50
rect 125 48 131 54
rect 125 46 127 48
rect 80 33 84 36
rect 70 32 84 33
rect 93 32 97 43
rect 101 38 107 46
rect 117 44 127 46
rect 117 42 131 44
rect 137 38 141 54
rect 101 34 104 38
rect 108 34 115 38
rect 119 34 120 38
rect 124 34 141 38
rect 74 28 84 32
rect 70 27 84 28
rect 44 18 53 22
rect 57 18 58 22
rect 36 12 40 18
rect 63 17 67 18
rect 73 22 77 23
rect 80 22 84 27
rect 87 31 97 32
rect 91 30 97 31
rect 91 29 122 30
rect 91 27 117 29
rect 87 26 117 27
rect 116 25 117 26
rect 121 25 122 29
rect 127 29 131 30
rect 80 18 90 22
rect 94 18 95 22
rect 106 18 107 22
rect 111 18 112 22
rect 73 12 77 18
rect 106 12 112 18
rect 127 12 131 25
rect 137 29 141 34
rect 137 24 141 25
rect -137 8 -131 12
rect -127 8 -64 12
rect -60 8 -36 12
rect -32 8 123 12
rect 127 8 134 12
rect 138 8 150 12
rect -137 4 150 8
<< ntransistor >>
rect -126 19 -124 30
rect -116 13 -114 30
rect -96 16 -94 30
rect -86 16 -84 30
rect -76 11 -74 30
rect -69 11 -67 30
rect -57 11 -55 30
rect -50 11 -48 30
rect -20 16 -18 30
rect -10 16 -8 30
rect 13 14 15 28
rect 31 23 33 30
rect 123 24 125 30
rect 42 17 44 23
rect 49 17 51 23
rect 59 17 61 23
rect 69 17 71 23
rect 79 17 81 23
rect 86 17 88 23
rect 96 17 98 23
rect 103 17 105 23
rect 133 23 135 30
<< ptransistor >>
rect -115 42 -113 70
rect -105 42 -103 70
rect -90 42 -88 70
rect -80 42 -78 70
rect -70 42 -68 55
rect -60 42 -58 55
rect -50 42 -48 70
rect -40 42 -38 70
rect -30 42 -28 70
rect -20 42 -18 70
rect -10 42 -8 70
rect 13 42 15 70
rect 23 42 25 56
rect 42 52 44 58
rect 49 52 51 58
rect 59 52 61 64
rect 69 52 71 64
rect 79 58 81 64
rect 86 58 88 64
rect 96 51 98 64
rect 103 51 105 64
rect 113 51 115 62
rect 133 53 135 63
<< polycontact >>
rect -63 59 -59 63
rect -125 34 -121 38
rect -79 34 -75 38
rect -49 34 -45 38
rect -33 34 -29 38
rect -13 34 -9 38
rect 14 33 18 37
rect 33 34 37 38
rect 50 43 54 47
rect 76 43 80 47
rect 56 27 60 31
rect 70 28 74 32
rect 93 43 97 47
rect 127 44 131 48
rect 87 27 91 31
rect 104 34 108 38
rect 120 34 124 38
<< ndcontact >>
rect -132 20 -128 24
rect -122 25 -118 29
rect -112 14 -108 18
rect -102 25 -98 29
rect -102 18 -98 22
rect -92 25 -88 29
rect -82 25 -78 29
rect -82 18 -78 22
rect -64 8 -60 12
rect -46 18 -42 22
rect -26 17 -22 21
rect -16 25 -12 29
rect -16 18 -12 22
rect 7 23 11 27
rect -6 17 -2 21
rect 25 25 29 29
rect 117 25 121 29
rect 127 25 131 29
rect 17 15 21 19
rect 36 18 40 22
rect 53 18 57 22
rect 63 18 67 22
rect 73 18 77 22
rect 90 18 94 22
rect 107 18 111 22
rect 137 25 141 29
<< pdcontact >>
rect -121 65 -117 69
rect -121 58 -117 62
rect -111 50 -107 54
rect -111 43 -107 47
rect -99 65 -95 69
rect -99 58 -95 62
rect -86 58 -82 62
rect -86 51 -82 55
rect -76 50 -72 54
rect -76 43 -72 47
rect -66 43 -62 47
rect -56 50 -52 54
rect -46 59 -42 63
rect -46 43 -42 47
rect -36 58 -32 62
rect -36 51 -32 55
rect -26 50 -22 54
rect -26 43 -22 47
rect -16 65 -12 69
rect -16 58 -12 62
rect -6 50 -2 54
rect -6 43 -2 47
rect 7 50 11 54
rect 7 43 11 47
rect 17 65 21 69
rect 17 51 21 55
rect 35 53 39 57
rect 53 53 57 57
rect 63 53 67 57
rect 73 59 77 63
rect 90 59 94 63
rect 27 43 31 47
rect 107 57 111 61
rect 127 58 131 62
rect 117 52 121 56
rect 137 54 141 58
<< psubstratepcontact >>
rect -131 8 -127 12
rect -36 8 -32 12
rect 123 8 127 12
rect 134 8 138 12
<< nsubstratencontact >>
rect -131 68 -127 72
rect -66 68 -62 72
rect 31 68 35 72
rect 41 68 45 72
rect 122 68 126 72
<< psubstratepdiff >>
rect -132 12 -126 13
rect -132 8 -131 12
rect -127 8 -126 12
rect -132 7 -126 8
rect -37 12 -31 28
rect -37 8 -36 12
rect -32 8 -31 12
rect -37 7 -31 8
rect 116 12 145 13
rect 116 8 123 12
rect 127 8 134 12
rect 138 8 145 12
rect 116 7 145 8
<< nsubstratendiff >>
rect -132 72 -126 73
rect -132 68 -131 72
rect -127 68 -126 72
rect -67 72 -61 73
rect -132 44 -126 68
rect -67 68 -66 72
rect -62 68 -61 72
rect 26 72 50 73
rect -67 67 -61 68
rect 26 68 31 72
rect 35 68 41 72
rect 45 68 50 72
rect 26 67 50 68
rect 121 72 127 73
rect 121 68 122 72
rect 126 68 127 72
rect 121 67 127 68
<< labels >>
rlabel polycontact 16 35 16 35 6 zn
rlabel polycontact 34 36 34 36 6 n4
rlabel polycontact 58 29 58 29 6 ci
rlabel polycontact 52 45 52 45 6 ci
rlabel polycontact 72 30 72 30 6 n1
rlabel polycontact 89 29 89 29 6 ci
rlabel polycontact 95 45 95 45 6 ci
rlabel polycontact 78 45 78 45 6 n2
rlabel polycontact 122 36 122 36 6 cn
rlabel metal1 21 35 21 35 6 zn
rlabel metal1 27 35 27 35 6 zn
rlabel metal1 51 20 51 20 6 n4
rlabel polycontact 57 29 57 29 6 ci
rlabel metal1 40 36 40 36 6 n4
rlabel polycontact 53 45 53 45 6 ci
rlabel metal1 50 55 50 55 6 n4
rlabel metal1 76 8 76 8 6 vss
rlabel metal1 77 30 77 30 6 n1
rlabel metal1 72 45 72 45 6 n2
rlabel metal1 65 37 65 37 6 n2
rlabel metal1 76 72 76 72 6 vdd
rlabel metal1 87 20 87 20 6 n1
rlabel metal1 112 36 112 36 6 d
rlabel metal1 104 40 104 40 6 d
rlabel metal1 95 40 95 40 6 ci
rlabel metal1 90 61 90 61 6 n1
rlabel metal1 104 28 104 28 6 ci
rlabel metal1 130 36 130 36 6 cn
rlabel metal1 120 44 120 44 6 cp
rlabel metal1 128 48 128 48 6 cp
rlabel metal1 139 41 139 41 6 cn
rlabel pdcontact 119 53 119 53 6 ci
rlabel polycontact -47 36 -47 36 6 an
rlabel polycontact -61 61 -61 61 6 bn
rlabel polycontact -31 36 -31 36 6 bn
rlabel polycontact -123 36 -123 36 6 b
rlabel metal1 -131 40 -131 40 6 b
rlabel metal1 -91 20 -91 20 6 z
rlabel metal1 -116 27 -116 27 6 bn
rlabel ndcontact -99 28 -99 28 6 z
rlabel metal1 -90 31 -90 31 6 an
rlabel metal1 -91 44 -91 44 6 z
rlabel metal1 -110 39 -110 39 6 bn
rlabel metal1 -84 56 -84 56 6 bn
rlabel metal1 -67 8 -67 8 6 vss
rlabel metal1 -59 20 -59 20 6 z
rlabel metal1 -67 20 -67 20 6 z
rlabel metal1 -75 20 -75 20 6 z
rlabel metal1 -83 20 -83 20 6 z
rlabel metal1 -83 44 -83 44 6 z
rlabel pdcontact -75 44 -75 44 6 z
rlabel metal1 -64 40 -64 40 6 an
rlabel metal1 -59 52 -59 52 6 z
rlabel metal1 -67 52 -67 52 6 z
rlabel metal1 -67 72 -67 72 6 vdd
rlabel ndcontact -43 20 -43 20 6 z
rlabel metal1 -51 20 -51 20 6 z
rlabel metal1 -34 40 -34 40 6 bn
rlabel metal1 -68 36 -68 36 6 an
rlabel pdcontact -44 44 -44 44 6 bn
rlabel metal1 -51 52 -51 52 6 z
rlabel metal1 -35 56 -35 56 6 z
rlabel metal1 -43 52 -43 52 6 z
rlabel metal1 -64 61 -64 61 6 bn
rlabel metal1 -14 23 -14 23 6 an
rlabel polycontact -11 36 -11 36 6 a
rlabel metal1 -4 49 -4 49 6 an
rlabel metal1 -14 45 -14 45 6 an
rlabel metal1 -25 49 -25 49 6 an
rlabel metal1 -3 32 -3 32 6 a
rlabel metal1 8 40 8 40 1 q
rlabel metal1 16 44 16 44 1 q
<< end >>
