* Tue Aug 10 11:21:07 CEST 2004
.subckt nd3_x4 a b c vdd vss z 
*SPICE circuit <nd3_x4> from XCircuit v3.10

m1 n1 a vss vss n w=66u l=2.3636u ad='66u*5u+12p' as='66u*5u+12p' pd='66u*2+14u' ps='66u*2+14u'
m2 n2 b n1 vss n w=66u l=2.3636u ad='66u*5u+12p' as='66u*5u+12p' pd='66u*2+14u' ps='66u*2+14u'
m3 z c n2 vss n w=66u l=2.3636u ad='66u*5u+12p' as='66u*5u+12p' pd='66u*2+14u' ps='66u*2+14u'
m4 z a vdd vdd p w=66u l=2.3636u ad='66u*5u+12p' as='66u*5u+12p' pd='66u*2+14u' ps='66u*2+14u'
m5 z b vdd vdd p w=66u l=2.3636u ad='66u*5u+12p' as='66u*5u+12p' pd='66u*2+14u' ps='66u*2+14u'
m6 z c vdd vdd p w=66u l=2.3636u ad='66u*5u+12p' as='66u*5u+12p' pd='66u*2+14u' ps='66u*2+14u'
.ends
