* Spice description of aoi22_x05
* Spice driver version 134999461
* Date 31/05/2007 at 21:32:39
* vxlib 0.13um values
.subckt aoi22_x05 a1 a2 b1 b2 vdd vss z
M1  sig5  b1    z     vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M2  vdd   a1    sig5  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M3  z     b2    sig5  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M4  sig5  a2    vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M5  n2    b1    vss   vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M6  vss   a1    sig3  vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M7  z     b2    n2    vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M8  sig3  a2    z     vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
C10 a1    vss   0.634f
C7  a2    vss   0.679f
C9  b1    vss   0.764f
C8  b2    vss   0.693f
C5  sig5  vss   0.574f
C4  z     vss   1.003f
.ends
