* Thu Jan 11 12:55:49 CET 2007
.subckt nd2av0x2 a b vdd vss z
*SPICE circuit <nd2av0x2> from XCircuit v3.20

m1 an a vss vss n w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m2 n1 b vss vss n w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m3 an a vdd vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m4 z b vdd vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m5 z an n1 vss n w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m6 z an vdd vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
.ends
