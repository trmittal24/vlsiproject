* Sun Apr  2 21:55:59 CEST 2006
.subckt nd2v3x05 a b vdd vss z 
*SPICE circuit <nd2v3x05> from XCircuit v3.20

m1 n1 a vss vss n w=17u l=2u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m2 z a vdd vdd p w=10u l=2u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m3 z b n1 vss n w=17u l=2u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m4 z b vdd vdd p w=10u l=2u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
.ends
