* Spice description of vddtie
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:11
*
.subckt vddtie vdd vss z 
C3  vdd   vss   0.477f
C1  z     vss   1.920f
.ends
