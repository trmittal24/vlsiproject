* Mon Aug 16 14:11:02 CEST 2004
.subckt or4v0x2 a b c d vdd vss z 
*SPICE circuit <or4v0x2> from XCircuit v3.10

m1 zn a vss vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m2 zn b vss vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m3 zn c vss vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m4 zn d n3 vdd p w=48u l=2u ad='48u*5u+12p' as='48u*5u+12p' pd='48u*2+14u' ps='48u*2+14u'
m5 n3 c n2 vdd p w=48u l=2u ad='48u*5u+12p' as='48u*5u+12p' pd='48u*2+14u' ps='48u*2+14u'
m6 n2 b n1 vdd p w=48u l=2u ad='48u*5u+12p' as='48u*5u+12p' pd='48u*2+14u' ps='48u*2+14u'
m7 n1 a vdd vdd p w=48u l=2u ad='48u*5u+12p' as='48u*5u+12p' pd='48u*2+14u' ps='48u*2+14u'
m8 z zn vss vss n w=14u l=2u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m9 z zn vdd vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m10 zn d vss vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
.ends
