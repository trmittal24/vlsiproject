magic
tech scmos
timestamp 1523164968
<< metal1 >>
rect 70 68 77 76
rect 141 68 150 76
rect -30 34 -27 38
rect 226 35 229 39
rect -30 24 -27 28
rect -30 14 -27 18
rect -6 8 4 12
rect -30 4 -27 8
rect -6 5 7 8
rect 70 5 77 12
rect 142 5 151 12
rect -6 4 214 5
rect -54 -7 -27 -3
rect -30 -17 -27 -13
rect -30 -27 -27 -23
rect -38 -37 -27 -33
rect -27 -58 -23 -45
rect -18 -57 -14 4
rect 2 -5 214 4
rect 70 -12 214 -5
rect 225 -40 229 -36
rect -4 -73 4 -68
rect -4 -75 5 -73
rect 70 -75 76 -68
rect 141 -75 147 -68
rect -4 -76 214 -75
rect 2 -92 214 -76
rect 225 -122 229 -118
rect -3 -156 5 -148
rect 68 -156 185 -148
<< metal2 >>
rect -26 45 61 46
rect -26 43 65 45
rect 71 44 133 47
rect 71 43 137 44
rect 141 44 205 47
rect 141 43 209 44
rect -26 38 -23 43
rect 71 38 74 43
rect 141 38 145 43
rect 10 34 74 38
rect 82 34 145 38
rect 154 35 222 39
rect -50 24 -27 28
rect -4 26 51 27
rect -4 24 55 26
rect -58 -147 -54 -7
rect -50 -49 -46 24
rect -4 18 -1 24
rect -42 14 -27 18
rect -23 14 -1 18
rect -42 -33 -38 14
rect -23 4 -18 8
rect 124 -3 128 26
rect -23 -7 128 -3
rect -34 -17 -27 -13
rect -34 -42 -31 -17
rect 15 -22 35 -18
rect 15 -23 18 -22
rect -23 -27 18 -23
rect 31 -23 35 -22
rect 82 -20 106 -17
rect 82 -23 85 -20
rect 31 -27 85 -23
rect 103 -23 106 -20
rect 197 -23 201 26
rect 103 -26 201 -23
rect 103 -27 160 -26
rect 164 -27 201 -26
rect 23 -33 26 -30
rect -23 -37 26 -33
rect 94 -34 98 -30
rect 66 -38 98 -34
rect -34 -45 -27 -42
rect 138 -42 146 -38
rect -23 -44 12 -42
rect 143 -43 146 -42
rect -23 -45 7 -44
rect 80 -49 84 -48
rect 143 -45 155 -43
rect 143 -49 151 -45
rect -50 -53 0 -49
rect -4 -54 0 -53
rect 17 -53 84 -49
rect 17 -54 21 -53
rect -27 -131 -23 -62
rect -4 -58 21 -54
rect -18 -80 -14 -61
rect -18 -84 65 -80
rect 62 -111 65 -84
rect 127 -115 133 -111
rect 197 -112 201 -27
rect 210 -40 221 -36
rect 197 -115 205 -112
rect 69 -119 92 -118
rect 127 -119 130 -115
rect 10 -121 130 -119
rect 10 -122 72 -121
rect 89 -122 130 -121
rect 154 -122 221 -119
rect 82 -129 186 -126
rect 182 -131 186 -129
rect -27 -135 53 -131
rect 182 -134 197 -131
rect 126 -147 130 -137
rect -58 -151 130 -147
<< m2contact >>
rect 61 45 65 49
rect 133 44 137 48
rect 205 44 209 48
rect -27 34 -23 38
rect 6 34 10 38
rect 78 34 82 38
rect 150 35 154 39
rect 222 35 226 39
rect -27 24 -23 28
rect 51 26 55 30
rect 124 26 128 30
rect 197 26 201 30
rect -27 14 -23 18
rect -27 4 -23 8
rect -18 4 -14 8
rect -58 -7 -54 -3
rect -27 -7 -23 -3
rect -27 -17 -23 -13
rect -27 -27 -23 -23
rect -42 -37 -38 -33
rect -27 -37 -23 -33
rect -27 -45 -23 -41
rect -27 -62 -23 -58
rect 23 -30 27 -26
rect 94 -30 98 -26
rect 160 -30 164 -26
rect 62 -38 66 -34
rect 134 -42 138 -38
rect 206 -40 210 -36
rect 221 -40 225 -36
rect 7 -49 12 -44
rect 80 -48 84 -44
rect 151 -49 155 -45
rect -18 -61 -14 -57
rect 61 -115 65 -111
rect 133 -115 137 -111
rect 205 -115 209 -111
rect 6 -123 10 -119
rect 150 -122 154 -118
rect 221 -122 225 -118
rect 78 -129 82 -125
rect 53 -135 57 -131
rect 126 -137 130 -133
rect 197 -134 201 -130
use or2v0x3  or2v0x3_0
timestamp 1521380365
transform 1 0 4 0 1 4
box -4 -4 68 76
use or2v0x3  or2v0x3_1
timestamp 1521380365
transform 1 0 76 0 1 4
box -4 -4 68 76
use or2v0x3  or2v0x3_2
timestamp 1521380365
transform 1 0 148 0 1 4
box -4 -4 68 76
use or2v0x3  or2v0x3_3
timestamp 1521380365
transform -1 0 68 0 -1 -4
box -4 -4 68 76
use or2v0x3  or2v0x3_4
timestamp 1521380365
transform -1 0 140 0 -1 -4
box -4 -4 68 76
use or2v0x3  or2v0x3_5
timestamp 1521380365
transform -1 0 212 0 -1 -4
box -4 -4 68 76
use or2v0x3  or2v0x3_6
timestamp 1521380365
transform 1 0 4 0 1 -156
box -4 -4 68 76
use or2v0x3  or2v0x3_7
timestamp 1521380365
transform 1 0 76 0 1 -156
box -4 -4 68 76
use or2v0x3  or2v0x3_8
timestamp 1521380365
transform 1 0 148 0 1 -156
box -4 -4 68 76
<< labels >>
rlabel metal1 -28 36 -28 36 3 d0
rlabel metal1 -29 16 -29 16 3 d2
rlabel metal1 -29 26 -29 26 3 d1
rlabel metal1 -29 6 -29 6 3 d3
rlabel metal1 -29 -5 -29 -5 3 d4
rlabel metal1 -29 -15 -29 -15 3 d5
rlabel metal1 -29 -25 -29 -25 3 d6
rlabel metal1 -3 8 -3 8 1 gnd
rlabel metal1 -2 72 -2 72 1 vdd
rlabel metal1 228 37 228 37 7 b0
rlabel metal1 227 -38 227 -38 7 b1
rlabel metal1 227 -120 227 -120 7 b2
rlabel metal1 -2 -72 -2 -72 1 vdd
rlabel metal1 -1 -153 -1 -153 1 gnd
<< end >>
