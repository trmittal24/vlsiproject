magic
tech scmos
timestamp 1521461618
<< pwell >>
rect 35 7 78 12
rect 2 -7 78 7
rect 35 -12 78 -7
<< polysilicon >>
rect 183 77 187 79
rect 183 72 185 77
<< metal1 >>
rect 182 79 183 83
rect -15 71 7 76
rect -15 -73 -11 71
rect 34 68 46 76
rect 77 68 83 76
rect 155 68 165 76
rect 205 68 215 76
rect 150 34 152 38
rect 242 34 244 38
rect -6 -7 -2 10
rect 35 7 88 12
rect 133 7 214 12
rect 2 2 254 7
rect 6 -2 254 2
rect 2 -5 254 -2
rect 2 -7 78 -5
rect 35 -12 78 -7
rect 84 -12 254 -5
rect 228 -30 237 -26
rect 50 -38 55 -34
rect 79 -38 103 -34
rect 142 -38 152 -34
rect 127 -46 137 -43
rect 31 -54 37 -50
rect 41 -54 48 -50
rect 93 -51 98 -47
rect 34 -72 46 -68
rect 84 -72 93 -68
rect 131 -72 141 -68
rect 213 -72 220 -68
rect 2 -73 270 -72
rect -15 -76 270 -73
rect -15 -230 -11 -76
rect 2 -91 270 -76
rect 2 -92 58 -91
rect 238 -92 270 -91
rect 73 -117 74 -113
rect 31 -126 36 -122
rect 1 -150 58 -148
rect 1 -160 227 -150
rect 5 -164 227 -160
rect 1 -172 227 -164
rect -15 -236 7 -230
rect 55 -236 177 -228
<< metal2 >>
rect -6 79 178 82
rect -6 14 -3 79
rect 163 47 200 50
rect 157 38 160 44
rect 252 42 256 45
rect 7 16 10 32
rect 46 21 49 32
rect 85 32 86 35
rect 125 32 139 35
rect 156 35 160 38
rect 136 30 139 32
rect 211 32 214 36
rect 136 27 159 30
rect 46 18 141 21
rect 7 13 40 16
rect -22 -1 2 2
rect -22 -161 -19 -1
rect -6 -111 -3 -11
rect 37 -35 40 13
rect 142 0 145 18
rect 142 -3 149 0
rect 21 -38 46 -35
rect 21 -73 24 -38
rect 89 -47 92 -29
rect 146 -34 149 -3
rect 156 -26 159 27
rect 166 26 169 31
rect 245 26 248 34
rect 166 23 248 26
rect 253 7 256 42
rect 206 4 256 7
rect 130 -37 138 -34
rect 38 -60 41 -54
rect 130 -60 133 -37
rect 146 -36 174 -34
rect 146 -37 178 -36
rect 206 -35 209 4
rect 222 -30 224 -26
rect 220 -42 228 -39
rect 38 -63 133 -60
rect 138 -62 141 -46
rect 220 -62 223 -42
rect 138 -65 223 -62
rect 21 -76 43 -73
rect 40 -101 43 -76
rect 40 -104 77 -101
rect 40 -110 43 -104
rect -6 -114 24 -111
rect 74 -113 77 -104
rect 104 -105 106 -101
rect 104 -111 107 -105
rect 21 -122 24 -114
rect 100 -114 107 -111
rect 21 -125 36 -122
rect -22 -164 1 -161
<< metal3 >>
rect 156 50 164 51
rect 156 44 157 50
rect 163 44 164 50
rect 156 43 164 44
rect 77 35 86 36
rect 77 29 79 35
rect 85 29 86 35
rect 77 1 86 29
rect 77 -7 92 1
rect 156 -5 162 43
rect 203 37 212 39
rect 203 31 205 37
rect 211 31 212 37
rect 203 29 213 31
rect 204 16 213 29
rect 204 10 220 16
rect 86 -22 92 -7
rect 130 -11 162 -5
rect 84 -23 94 -22
rect 84 -29 86 -23
rect 92 -29 94 -23
rect 84 -31 94 -29
rect 130 -73 137 -11
rect 214 -24 220 10
rect 214 -26 223 -24
rect 214 -32 216 -26
rect 222 -32 223 -26
rect 214 -34 223 -32
rect 105 -80 137 -73
rect 105 -99 113 -80
rect 105 -105 106 -99
rect 112 -105 113 -99
rect 105 -106 113 -105
<< polycontact >>
rect 183 79 187 83
<< m2contact >>
rect 178 79 182 83
rect 200 46 204 50
rect 248 42 252 46
rect 6 32 10 36
rect 46 32 50 36
rect 86 32 90 36
rect 121 32 125 36
rect 152 34 156 38
rect 166 31 170 35
rect 214 32 218 36
rect 244 34 248 38
rect 141 18 145 22
rect -6 10 -2 14
rect 2 -2 6 2
rect -6 -11 -2 -7
rect 156 -30 160 -26
rect 224 -30 228 -26
rect 46 -38 50 -34
rect 138 -38 142 -34
rect 174 -36 178 -32
rect 206 -39 210 -35
rect 228 -42 232 -38
rect 137 -46 141 -42
rect 37 -54 41 -50
rect 89 -51 93 -47
rect 40 -114 44 -110
rect 74 -117 78 -113
rect 96 -115 100 -111
rect 36 -126 40 -122
rect 1 -164 5 -160
<< m3contact >>
rect 157 44 163 50
rect 79 29 85 35
rect 205 31 211 37
rect 86 -29 92 -23
rect 216 -32 222 -26
rect 106 -105 112 -99
use ../pharosc_8.4/magic/cells/vsclib/iv1v0x4  iv1v0x4_0
timestamp 1521461618
transform 1 0 4 0 1 4
box -4 -4 36 76
use ../pharosc_8.4/magic/cells/vsclib/iv1v0x4  iv1v0x4_1
timestamp 1521461618
transform 1 0 44 0 1 4
box -4 -4 36 76
use ../pharosc_8.4/magic/cells/vsclib/or3v0x2  or3v0x2_0
timestamp 1521461618
transform 1 0 84 0 1 4
box -4 -4 76 76
use ../pharosc_8.4/magic/cells/vsclib/an2v0x2  an2v0x2_2
timestamp 1521461618
transform 1 0 164 0 1 4
box -4 -4 44 76
use ../pharosc_8.4/magic/cells/vsclib/an2v0x2  an2v0x2_3
timestamp 1521461618
transform 1 0 212 0 1 4
box -4 -4 44 76
use ../pharosc_8.4/magic/cells/vsclib/iv1v0x4  iv1v0x4_2
timestamp 1521461618
transform -1 0 36 0 -1 -4
box -4 -4 36 76
use ../pharosc_8.4/magic/cells/vsclib/an2v0x2  an2v0x2_0
timestamp 1521461618
transform -1 0 84 0 -1 -4
box -4 -4 44 76
use ../pharosc_8.4/magic/cells/vsclib/an2v0x2  an2v0x2_1
timestamp 1521461618
transform -1 0 132 0 -1 -4
box -4 -4 44 76
use ../pharosc_8.4/magic/cells/vsclib/or3v0x2  or3v0x2_1
timestamp 1521461618
transform -1 0 212 0 -1 -4
box -4 -4 76 76
use ../pharosc_8.4/magic/cells/vsclib/nr2v0x2  nr2v0x2_0
timestamp 1521461618
transform -1 0 268 0 -1 -4
box -4 -4 52 76
use ../pharosc_8.4/magic/cells/vsclib/an2v0x2  an2v0x2_4
timestamp 1521461618
transform 1 0 4 0 1 -156
box -4 -4 44 76
use ../pharosc_8.4/magic/cells/vsclib/an3v0x2  an3v0x2_0
timestamp 1521461618
transform 1 0 52 0 1 -156
box -4 -4 60 76
use ../pharosc_8.4/magic/cells/vsclib/an3v0x2  an3v0x2_3
timestamp 1521461618
transform 1 0 116 0 1 -156
box -4 -4 60 76
use ../pharosc_8.4/magic/cells/vsclib/nr2v0x2  nr2v0x2_1
timestamp 1521461618
transform 1 0 180 0 1 -156
box -4 -4 52 76
use ../pharosc_8.4/magic/cells/vsclib/an3v0x2  an3v0x2_2
timestamp 1521461618
transform -1 0 60 0 -1 -164
box -4 -4 60 76
use ../pharosc_8.4/magic/cells/vsclib/nr3v0x2  nr3v0x2_0
timestamp 1521461618
transform -1 0 156 0 -1 -164
box -4 -4 92 76
use ../pharosc_8.4/magic/cells/vsclib/an3v0x2  an3v0x2_1
timestamp 1521461618
transform -1 0 220 0 -1 -164
box -4 -4 60 76
<< end >>
