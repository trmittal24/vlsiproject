* Sat Aug 27 22:09:57 CEST 2005
.subckt iv1v4x1 a vdd vss z 
*SPICE circuit <iv1v4x1> from XCircuit v3.20

m1 z a vss vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m2 z a vdd vdd p w=24u l=2.3636u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
.ends
