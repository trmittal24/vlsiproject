* SPICE3 file created from subcomp.ext - technology: scmos
.include t14y_tsmc_025_level3.txt

M1000 comp_0_nd3v0x2_0_z comp_0_nr3v0x2_0_z totdiff3_0_mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=14u l=2u
+  ad=392p pd=120u as=31188p ps=11196u
M1001 totdiff3_0_mux_0_vdd comp_0_nr3v0x2_0_z comp_0_nd3v0x2_0_z comp_0_an3v0x2_2_w_n4_32# pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1002 comp_0_nd3v0x2_0_z comp_0_nd3v0x2_0_c totdiff3_0_mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1003 totdiff3_0_mux_0_vdd comp_0_nd3v0x2_0_a comp_0_nd3v0x2_0_z comp_0_an3v0x2_2_w_n4_32# pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1004 comp_0_nd3v0x2_0_a_14_12# comp_0_nd3v0x2_0_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=70p pd=38u as=21022p ps=7450u
M1005 comp_0_nd3v0x2_0_a_21_12# comp_0_nr3v0x2_0_z comp_0_nd3v0x2_0_a_14_12# totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=70p pd=38u as=0p ps=0u
M1006 comp_0_nd3v0x2_0_z comp_0_nd3v0x2_0_c comp_0_nd3v0x2_0_a_21_12# totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=112p pd=44u as=0p ps=0u
M1007 comp_0_nd3v0x2_0_a_38_12# comp_0_nd3v0x2_0_c comp_0_nd3v0x2_0_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=70p pd=38u as=0p ps=0u
M1008 comp_0_nd3v0x2_0_a_45_12# comp_0_nr3v0x2_0_z comp_0_nd3v0x2_0_a_38_12# totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=70p pd=38u as=0p ps=0u
M1009 totdiff3_0_mux_0_gnd comp_0_nd3v0x2_0_a comp_0_nd3v0x2_0_a_45_12# totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1010 totdiff3_0_mux_0_vdd comp_0_an3v0x2_1_zn comp_0_nr2v0x2_1_a comp_0_an3v0x2_2_w_n4_32# pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1011 comp_0_an3v0x2_1_zn comp_0_an3v0x2_1_a totdiff3_0_mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=17u l=2u
+  ad=233p pd=98u as=0p ps=0u
M1012 totdiff3_0_mux_0_vdd comp_0_an3v0x2_2_b comp_0_an3v0x2_1_zn comp_0_an3v0x2_2_w_n4_32# pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1013 comp_0_an3v0x2_1_zn comp_0_an3v0x2_2_c totdiff3_0_mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1014 totdiff3_0_mux_0_gnd comp_0_an3v0x2_1_zn comp_0_nr2v0x2_1_a totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=82p ps=42u
M1015 comp_0_an3v0x2_1_a_24_8# comp_0_an3v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1016 comp_0_an3v0x2_1_a_31_8# comp_0_an3v0x2_2_b comp_0_an3v0x2_1_a_24_8# totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1017 comp_0_an3v0x2_1_zn comp_0_an3v0x2_2_c comp_0_an3v0x2_1_a_31_8# totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=97p pd=48u as=0p ps=0u
M1018 comp_0_nr3v0x2_0_a_13_39# comp_0_an3v0x2_2_z comp_0_nr3v0x2_0_z comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=135p pd=64u as=377p ps=138u
M1019 comp_0_nr3v0x2_0_a_20_39# comp_0_an3v0x2_0_z comp_0_nr3v0x2_0_a_13_39# comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1020 totdiff3_0_mux_0_vdd comp_0_nr3v0x2_0_a comp_0_nr3v0x2_0_a_20_39# comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1021 comp_0_nr3v0x2_0_a_37_39# comp_0_nr3v0x2_0_a totdiff3_0_mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1022 comp_0_nr3v0x2_0_a_44_39# comp_0_an3v0x2_0_z comp_0_nr3v0x2_0_a_37_39# comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1023 comp_0_nr3v0x2_0_z comp_0_an3v0x2_2_z comp_0_nr3v0x2_0_a_44_39# comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1024 comp_0_nr3v0x2_0_a_61_39# comp_0_an3v0x2_2_z comp_0_nr3v0x2_0_z comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1025 comp_0_nr3v0x2_0_a_68_39# comp_0_an3v0x2_0_z comp_0_nr3v0x2_0_a_61_39# comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1026 totdiff3_0_mux_0_vdd comp_0_nr3v0x2_0_a comp_0_nr3v0x2_0_a_68_39# comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1027 totdiff3_0_mux_0_gnd comp_0_an3v0x2_2_z comp_0_nr3v0x2_0_z totdiff3_0_mux_0_gnd nfet w=15u l=2u
+  ad=0p pd=0u as=207p ps=90u
M1028 comp_0_nr3v0x2_0_z comp_0_an3v0x2_0_z totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=15u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1029 totdiff3_0_mux_0_gnd comp_0_nr3v0x2_0_a comp_0_nr3v0x2_0_z totdiff3_0_mux_0_gnd nfet w=15u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1030 totdiff3_0_mux_0_vdd comp_0_an3v0x2_2_zn comp_0_an3v0x2_2_z comp_0_an3v0x2_2_w_n4_32# pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1031 comp_0_an3v0x2_2_zn comp_0_an3v0x2_2_a totdiff3_0_mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=17u l=2u
+  ad=233p pd=98u as=0p ps=0u
M1032 totdiff3_0_mux_0_vdd comp_0_an3v0x2_2_b comp_0_an3v0x2_2_zn comp_0_an3v0x2_2_w_n4_32# pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1033 comp_0_an3v0x2_2_zn comp_0_an3v0x2_2_c totdiff3_0_mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1034 totdiff3_0_mux_0_gnd comp_0_an3v0x2_2_zn comp_0_an3v0x2_2_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=82p ps=42u
M1035 comp_0_an3v0x2_2_a_24_8# comp_0_an3v0x2_2_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1036 comp_0_an3v0x2_2_a_31_8# comp_0_an3v0x2_2_b comp_0_an3v0x2_2_a_24_8# totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1037 comp_0_an3v0x2_2_zn comp_0_an3v0x2_2_c comp_0_an3v0x2_2_a_31_8# totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=97p pd=48u as=0p ps=0u
M1038 comp_0_nr2v0x2_1_a_11_39# comp_0_nr2v0x2_1_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1039 comp_0_nd3v0x2_0_c comp_0_an3v0x2_3_z comp_0_nr2v0x2_1_a_11_39# totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=216p pd=70u as=0p ps=0u
M1040 comp_0_nr2v0x2_1_a_28_39# comp_0_an3v0x2_3_z comp_0_nd3v0x2_0_c totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1041 totdiff3_0_mux_0_vdd comp_0_nr2v0x2_1_a comp_0_nr2v0x2_1_a_28_39# totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1042 comp_0_nd3v0x2_0_c comp_0_nr2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=15u l=2u
+  ad=120p pd=46u as=0p ps=0u
M1043 totdiff3_0_mux_0_gnd comp_0_an3v0x2_3_z comp_0_nd3v0x2_0_c totdiff3_0_mux_0_gnd nfet w=15u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1044 totdiff3_0_mux_0_vdd comp_0_an3v0x2_3_zn comp_0_an3v0x2_3_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1045 comp_0_an3v0x2_3_zn comp_0_an2v0x2_0_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=17u l=2u
+  ad=233p pd=98u as=0p ps=0u
M1046 totdiff3_0_mux_0_vdd comp_0_an3v0x2_0_b comp_0_an3v0x2_3_zn totdiff3_0_mux_0_vdd pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1047 comp_0_an3v0x2_3_zn comp_0_an3v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1048 totdiff3_0_mux_0_gnd comp_0_an3v0x2_3_zn comp_0_an3v0x2_3_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=82p ps=42u
M1049 comp_0_an3v0x2_3_a_24_8# comp_0_an2v0x2_0_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1050 comp_0_an3v0x2_3_a_31_8# comp_0_an3v0x2_0_b comp_0_an3v0x2_3_a_24_8# totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1051 comp_0_an3v0x2_3_zn comp_0_an3v0x2_2_a comp_0_an3v0x2_3_a_31_8# totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=97p pd=48u as=0p ps=0u
M1052 totdiff3_0_mux_0_vdd comp_0_an3v0x2_0_zn comp_0_an3v0x2_0_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1053 comp_0_an3v0x2_0_zn comp_0_an3v0x2_1_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=17u l=2u
+  ad=233p pd=98u as=0p ps=0u
M1054 totdiff3_0_mux_0_vdd comp_0_an3v0x2_0_b comp_0_an3v0x2_0_zn totdiff3_0_mux_0_vdd pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1055 comp_0_an3v0x2_0_zn comp_0_an2v0x2_0_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1056 totdiff3_0_mux_0_gnd comp_0_an3v0x2_0_zn comp_0_an3v0x2_0_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=82p ps=42u
M1057 comp_0_an3v0x2_0_a_24_8# comp_0_an3v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1058 comp_0_an3v0x2_0_a_31_8# comp_0_an3v0x2_0_b comp_0_an3v0x2_0_a_24_8# totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1059 comp_0_an3v0x2_0_zn comp_0_an2v0x2_0_b comp_0_an3v0x2_0_a_31_8# totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=97p pd=48u as=0p ps=0u
M1060 totdiff3_0_mux_0_vdd comp_0_an2v0x2_0_zn comp_0_nr3v0x2_0_a totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1061 comp_0_an2v0x2_0_zn comp_0_an3v0x2_2_c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1062 totdiff3_0_mux_0_vdd comp_0_an2v0x2_0_b comp_0_an2v0x2_0_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1063 totdiff3_0_mux_0_gnd comp_0_an2v0x2_0_zn comp_0_nr3v0x2_0_a totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1064 comp_0_an2v0x2_0_a_24_13# comp_0_an3v0x2_2_c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1065 comp_0_an2v0x2_0_zn comp_0_an2v0x2_0_b comp_0_an2v0x2_0_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1066 comp_0_nr2v0x2_0_a_11_39# comp_0_an2v0x2_3_z totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1067 comp_0_nd3v0x2_0_a comp_0_an2v0x2_1_z comp_0_nr2v0x2_0_a_11_39# totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=216p pd=70u as=0p ps=0u
M1068 comp_0_nr2v0x2_0_a_28_39# comp_0_an2v0x2_1_z comp_0_nd3v0x2_0_a totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1069 totdiff3_0_mux_0_vdd comp_0_an2v0x2_3_z comp_0_nr2v0x2_0_a_28_39# totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1070 comp_0_nd3v0x2_0_a comp_0_an2v0x2_3_z totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=15u l=2u
+  ad=120p pd=46u as=0p ps=0u
M1071 totdiff3_0_mux_0_gnd comp_0_an2v0x2_1_z comp_0_nd3v0x2_0_a totdiff3_0_mux_0_gnd nfet w=15u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1072 totdiff3_0_mux_0_vdd comp_0_or3v0x2_1_zn comp_0_an2v0x2_3_b totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1073 comp_0_or3v0x2_1_a_24_38# comp_0_an3v0x2_2_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=22u l=2u
+  ad=110p pd=54u as=0p ps=0u
M1074 comp_0_or3v0x2_1_a_31_38# comp_0_an3v0x2_1_a comp_0_or3v0x2_1_a_24_38# totdiff3_0_mux_0_vdd pfet w=22u l=2u
+  ad=110p pd=54u as=0p ps=0u
M1075 comp_0_or3v0x2_1_zn comp_0_an3v0x2_2_a comp_0_or3v0x2_1_a_31_38# totdiff3_0_mux_0_vdd pfet w=22u l=2u
+  ad=167p pd=60u as=0p ps=0u
M1076 comp_0_or3v0x2_1_a_48_38# comp_0_an3v0x2_2_a comp_0_or3v0x2_1_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=95p pd=48u as=0p ps=0u
M1077 comp_0_or3v0x2_1_a_55_38# comp_0_an3v0x2_1_a comp_0_or3v0x2_1_a_48_38# totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=95p pd=48u as=0p ps=0u
M1078 totdiff3_0_mux_0_vdd comp_0_an3v0x2_2_b comp_0_or3v0x2_1_a_55_38# totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1079 totdiff3_0_mux_0_gnd comp_0_or3v0x2_1_zn comp_0_an2v0x2_3_b totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1080 comp_0_or3v0x2_1_zn comp_0_an3v0x2_2_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=8u l=2u
+  ad=116p pd=62u as=0p ps=0u
M1081 totdiff3_0_mux_0_gnd comp_0_an3v0x2_1_a comp_0_or3v0x2_1_zn totdiff3_0_mux_0_gnd nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1082 comp_0_or3v0x2_1_zn comp_0_an3v0x2_2_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1083 totdiff3_0_mux_0_vdd comp_0_an2v0x2_1_zn comp_0_an2v0x2_1_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1084 comp_0_an2v0x2_1_zn comp_0_an2v0x2_4_z totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1085 totdiff3_0_mux_0_vdd comp_0_an2v0x2_1_b comp_0_an2v0x2_1_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1086 totdiff3_0_mux_0_gnd comp_0_an2v0x2_1_zn comp_0_an2v0x2_1_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1087 comp_0_an2v0x2_1_a_24_13# comp_0_an2v0x2_4_z totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1088 comp_0_an2v0x2_1_zn comp_0_an2v0x2_1_b comp_0_an2v0x2_1_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1089 totdiff3_0_mux_0_vdd comp_0_an2v0x2_4_zn comp_0_an2v0x2_4_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1090 comp_0_an2v0x2_4_zn comp_0_an2v0x2_0_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1091 totdiff3_0_mux_0_vdd comp_0_an3v0x2_2_b comp_0_an2v0x2_4_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1092 totdiff3_0_mux_0_gnd comp_0_an2v0x2_4_zn comp_0_an2v0x2_4_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1093 comp_0_an2v0x2_4_a_24_13# comp_0_an2v0x2_0_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1094 comp_0_an2v0x2_4_zn comp_0_an3v0x2_2_b comp_0_an2v0x2_4_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1095 comp_0_an3v0x2_2_b comp_0_iv1v0x4_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1096 totdiff3_0_mux_0_vdd comp_0_iv1v0x4_2_a comp_0_an3v0x2_2_b totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1097 comp_0_an3v0x2_2_b comp_0_iv1v0x4_2_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=118p pd=50u as=0p ps=0u
M1098 totdiff3_0_mux_0_gnd comp_0_iv1v0x4_2_a comp_0_an3v0x2_2_b totdiff3_0_mux_0_gnd nfet w=11u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1099 totdiff3_0_mux_0_vdd comp_0_an2v0x2_3_zn comp_0_an2v0x2_3_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1100 comp_0_an2v0x2_3_zn comp_0_an2v0x2_2_z totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1101 totdiff3_0_mux_0_vdd comp_0_an2v0x2_3_b comp_0_an2v0x2_3_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1102 totdiff3_0_mux_0_gnd comp_0_an2v0x2_3_zn comp_0_an2v0x2_3_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1103 comp_0_an2v0x2_3_a_24_13# comp_0_an2v0x2_2_z totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1104 comp_0_an2v0x2_3_zn comp_0_an2v0x2_3_b comp_0_an2v0x2_3_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1105 totdiff3_0_mux_0_vdd comp_0_an2v0x2_2_zn comp_0_an2v0x2_2_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1106 comp_0_an2v0x2_2_zn comp_0_an3v0x2_2_c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1107 totdiff3_0_mux_0_vdd comp_0_an3v0x2_0_b comp_0_an2v0x2_2_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1108 totdiff3_0_mux_0_gnd comp_0_an2v0x2_2_zn comp_0_an2v0x2_2_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1109 comp_0_an2v0x2_2_a_24_13# comp_0_an3v0x2_2_c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1110 comp_0_an2v0x2_2_zn comp_0_an3v0x2_0_b comp_0_an2v0x2_2_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1111 totdiff3_0_mux_0_vdd comp_0_or3v0x2_0_zn comp_0_an2v0x2_1_b totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1112 comp_0_or3v0x2_0_a_24_38# comp_0_an3v0x2_0_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=22u l=2u
+  ad=110p pd=54u as=0p ps=0u
M1113 comp_0_or3v0x2_0_a_31_38# comp_0_an3v0x2_2_a comp_0_or3v0x2_0_a_24_38# totdiff3_0_mux_0_vdd pfet w=22u l=2u
+  ad=110p pd=54u as=0p ps=0u
M1114 comp_0_or3v0x2_0_zn comp_0_an3v0x2_1_a comp_0_or3v0x2_0_a_31_38# totdiff3_0_mux_0_vdd pfet w=22u l=2u
+  ad=167p pd=60u as=0p ps=0u
M1115 comp_0_or3v0x2_0_a_48_38# comp_0_an3v0x2_1_a comp_0_or3v0x2_0_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=95p pd=48u as=0p ps=0u
M1116 comp_0_or3v0x2_0_a_55_38# comp_0_an3v0x2_2_a comp_0_or3v0x2_0_a_48_38# totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=95p pd=48u as=0p ps=0u
M1117 totdiff3_0_mux_0_vdd comp_0_an3v0x2_0_b comp_0_or3v0x2_0_a_55_38# totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1118 totdiff3_0_mux_0_gnd comp_0_or3v0x2_0_zn comp_0_an2v0x2_1_b totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1119 comp_0_or3v0x2_0_zn comp_0_an3v0x2_0_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=8u l=2u
+  ad=116p pd=62u as=0p ps=0u
M1120 totdiff3_0_mux_0_gnd comp_0_an3v0x2_2_a comp_0_or3v0x2_0_zn totdiff3_0_mux_0_gnd nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1121 comp_0_or3v0x2_0_zn comp_0_an3v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1122 comp_0_an3v0x2_1_a comp_0_iv1v0x4_1_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1123 totdiff3_0_mux_0_vdd comp_0_iv1v0x4_1_a comp_0_an3v0x2_1_a totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1124 comp_0_an3v0x2_1_a comp_0_iv1v0x4_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=118p pd=50u as=0p ps=0u
M1125 totdiff3_0_mux_0_gnd comp_0_iv1v0x4_1_a comp_0_an3v0x2_1_a totdiff3_0_mux_0_gnd nfet w=11u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1126 comp_0_an2v0x2_0_b comp_0_iv1v0x4_0_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1127 totdiff3_0_mux_0_vdd comp_0_iv1v0x4_0_a comp_0_an2v0x2_0_b totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1128 comp_0_an2v0x2_0_b comp_0_iv1v0x4_0_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=17u l=2u
+  ad=118p pd=50u as=0p ps=0u
M1129 totdiff3_0_mux_0_gnd comp_0_iv1v0x4_0_a comp_0_an2v0x2_0_b totdiff3_0_mux_0_gnd nfet w=11u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1130 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_2_zn comp_0_iv1v0x4_0_a totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1131 totdiff3_1_mux_0_mxn2v0x1_2_a_21_50# totdiff3_1_mux_0_a2 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1132 totdiff3_1_mux_0_mxn2v0x1_2_zn totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_2_a_21_50# totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1133 totdiff3_1_mux_0_mxn2v0x1_2_a_38_50# totdiff3_1_mux_0_mxn2v0x1_2_sn totdiff3_1_mux_0_mxn2v0x1_2_zn totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1134 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_b2 totdiff3_1_mux_0_mxn2v0x1_2_a_38_50# totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1135 totdiff3_1_mux_0_mxn2v0x1_2_sn totdiff3_1_mux_0_s totdiff3_0_mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1136 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_2_zn comp_0_iv1v0x4_0_a totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1137 totdiff3_1_mux_0_mxn2v0x1_2_a_21_12# totdiff3_1_mux_0_a2 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1138 totdiff3_1_mux_0_mxn2v0x1_2_zn totdiff3_1_mux_0_mxn2v0x1_2_sn totdiff3_1_mux_0_mxn2v0x1_2_a_21_12# totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1139 totdiff3_1_mux_0_mxn2v0x1_2_a_38_12# totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_2_zn totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1140 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_b2 totdiff3_1_mux_0_mxn2v0x1_2_a_38_12# totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1141 totdiff3_1_mux_0_mxn2v0x1_2_sn totdiff3_1_mux_0_s totdiff3_0_mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1142 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_1_zn comp_0_iv1v0x4_2_a totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1143 totdiff3_1_mux_0_mxn2v0x1_1_a_21_50# totdiff3_1_mux_0_a1 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1144 totdiff3_1_mux_0_mxn2v0x1_1_zn totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_1_a_21_50# totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1145 totdiff3_1_mux_0_mxn2v0x1_1_a_38_50# totdiff3_1_mux_0_mxn2v0x1_1_sn totdiff3_1_mux_0_mxn2v0x1_1_zn totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1146 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_b1 totdiff3_1_mux_0_mxn2v0x1_1_a_38_50# totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1147 totdiff3_1_mux_0_mxn2v0x1_1_sn totdiff3_1_mux_0_s totdiff3_0_mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1148 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_1_zn comp_0_iv1v0x4_2_a totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1149 totdiff3_1_mux_0_mxn2v0x1_1_a_21_12# totdiff3_1_mux_0_a1 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1150 totdiff3_1_mux_0_mxn2v0x1_1_zn totdiff3_1_mux_0_mxn2v0x1_1_sn totdiff3_1_mux_0_mxn2v0x1_1_a_21_12# totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1151 totdiff3_1_mux_0_mxn2v0x1_1_a_38_12# totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_1_zn totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1152 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_b1 totdiff3_1_mux_0_mxn2v0x1_1_a_38_12# totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1153 totdiff3_1_mux_0_mxn2v0x1_1_sn totdiff3_1_mux_0_s totdiff3_0_mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1154 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_0_zn comp_0_iv1v0x4_1_a totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1155 totdiff3_1_mux_0_mxn2v0x1_0_a_21_50# totdiff3_1_mux_0_a0 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1156 totdiff3_1_mux_0_mxn2v0x1_0_zn totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_0_a_21_50# totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1157 totdiff3_1_mux_0_mxn2v0x1_0_a_38_50# totdiff3_1_mux_0_mxn2v0x1_0_sn totdiff3_1_mux_0_mxn2v0x1_0_zn totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1158 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_b0 totdiff3_1_mux_0_mxn2v0x1_0_a_38_50# totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1159 totdiff3_1_mux_0_mxn2v0x1_0_sn totdiff3_1_mux_0_s totdiff3_0_mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1160 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_0_zn comp_0_iv1v0x4_1_a totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1161 totdiff3_1_mux_0_mxn2v0x1_0_a_21_12# totdiff3_1_mux_0_a0 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1162 totdiff3_1_mux_0_mxn2v0x1_0_zn totdiff3_1_mux_0_mxn2v0x1_0_sn totdiff3_1_mux_0_mxn2v0x1_0_a_21_12# totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1163 totdiff3_1_mux_0_mxn2v0x1_0_a_38_12# totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_0_zn totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1164 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_b0 totdiff3_1_mux_0_mxn2v0x1_0_a_38_12# totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1165 totdiff3_1_mux_0_mxn2v0x1_0_sn totdiff3_1_mux_0_s totdiff3_0_mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1166 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_an2v0x2_2_zn totdiff3_1_diff2_2_an2v0x2_2_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1167 totdiff3_1_diff2_2_an2v0x2_2_zn totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1168 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_in_2c totdiff3_1_diff2_2_an2v0x2_2_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1169 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_an2v0x2_2_zn totdiff3_1_diff2_2_an2v0x2_2_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1170 totdiff3_1_diff2_2_an2v0x2_2_a_24_13# totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1171 totdiff3_1_diff2_2_an2v0x2_2_zn totdiff3_1_diff2_2_in_2c totdiff3_1_diff2_2_an2v0x2_2_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1172 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_mux_0_b2 totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1173 totdiff3_1_mux_0_b2 totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1174 totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_mux_0_b2 totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1175 totdiff3_1_mux_0_b2 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1176 totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_diff2_2_in_2c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1177 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_in_2c totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1178 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1179 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1180 totdiff3_1_diff2_2_xor2v2x2_0_a_13_13# totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1181 totdiff3_1_mux_0_b2 totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_diff2_2_xor2v2x2_0_a_13_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1182 totdiff3_1_diff2_2_xor2v2x2_0_a_30_13# totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_mux_0_b2 totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1183 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_diff2_2_xor2v2x2_0_a_30_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1184 totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_diff2_2_in_2c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1185 totdiff3_1_mux_0_b2 totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1186 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_diff2_2_in_2c totdiff3_1_mux_0_b2 totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1187 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1188 totdiff3_1_mux_0_s totdiff3_1_diff2_2_or2v0x3_0_zn totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1189 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_or2v0x3_0_zn totdiff3_1_mux_0_s totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1190 totdiff3_1_diff2_2_or2v0x3_0_a_31_39# totdiff3_1_diff2_2_an2v0x2_1_z totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1191 totdiff3_1_diff2_2_or2v0x3_0_zn totdiff3_1_diff2_2_an2v0x2_0_z totdiff3_1_diff2_2_or2v0x3_0_a_31_39# totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1192 totdiff3_1_diff2_2_or2v0x3_0_a_48_39# totdiff3_1_diff2_2_an2v0x2_0_z totdiff3_1_diff2_2_or2v0x3_0_zn totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1193 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_an2v0x2_1_z totdiff3_1_diff2_2_or2v0x3_0_a_48_39# totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1194 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_or2v0x3_0_zn totdiff3_1_mux_0_s totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1195 totdiff3_1_diff2_2_or2v0x3_0_zn totdiff3_1_diff2_2_an2v0x2_1_z totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1196 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_an2v0x2_0_z totdiff3_1_diff2_2_or2v0x3_0_zn totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1197 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_an2v0x2_1_zn totdiff3_1_diff2_2_an2v0x2_1_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1198 totdiff3_1_diff2_2_an2v0x2_1_zn totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1199 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_an2v0x2_1_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1200 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_an2v0x2_1_zn totdiff3_1_diff2_2_an2v0x2_1_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1201 totdiff3_1_diff2_2_an2v0x2_1_a_24_13# totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1202 totdiff3_1_diff2_2_an2v0x2_1_zn totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_an2v0x2_1_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1203 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_an2v0x2_0_zn totdiff3_1_diff2_2_an2v0x2_0_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1204 totdiff3_1_diff2_2_an2v0x2_0_zn totdiff3_1_diff2_2_in_c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1205 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_an2v0x2_0_b totdiff3_1_diff2_2_an2v0x2_0_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1206 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_an2v0x2_0_zn totdiff3_1_diff2_2_an2v0x2_0_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1207 totdiff3_1_diff2_2_an2v0x2_0_a_24_13# totdiff3_1_diff2_2_in_c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1208 totdiff3_1_diff2_2_an2v0x2_0_zn totdiff3_1_diff2_2_an2v0x2_0_b totdiff3_1_diff2_2_an2v0x2_0_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1209 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_xnr2v8x05_0_zn totdiff3_1_diff2_2_an2v0x2_0_b totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1210 totdiff3_1_diff2_2_xnr2v8x05_0_an totdiff3_1_diff2_2_in_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1211 totdiff3_1_diff2_2_xnr2v8x05_0_zn totdiff3_1_diff2_2_xnr2v8x05_0_bn totdiff3_1_diff2_2_xnr2v8x05_0_an totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1212 totdiff3_1_diff2_2_xnr2v8x05_0_ai totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_xnr2v8x05_0_zn totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1213 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_xnr2v8x05_0_an totdiff3_1_diff2_2_xnr2v8x05_0_ai totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1214 totdiff3_1_diff2_2_xnr2v8x05_0_bn totdiff3_1_diff2_2_in_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1215 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_xnr2v8x05_0_zn totdiff3_1_diff2_2_an2v0x2_0_b totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1216 totdiff3_1_diff2_2_xnr2v8x05_0_an totdiff3_1_diff2_2_in_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1217 totdiff3_1_diff2_2_xnr2v8x05_0_zn totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_xnr2v8x05_0_an totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1218 totdiff3_1_diff2_2_xnr2v8x05_0_ai totdiff3_1_diff2_2_xnr2v8x05_0_bn totdiff3_1_diff2_2_xnr2v8x05_0_zn totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1219 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_xnr2v8x05_0_an totdiff3_1_diff2_2_xnr2v8x05_0_ai totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1220 totdiff3_1_diff2_2_xnr2v8x05_0_bn totdiff3_1_diff2_2_in_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1221 totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_1_mux_0_a2 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1222 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1223 totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_1_mux_0_a2 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1224 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1225 totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_mux_0_a2 totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1226 totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1227 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_mux_0_a2 totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1228 totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1229 totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_diff2_2_in_c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1230 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_in_c totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_0_mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1231 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1232 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1233 totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_1_diff2_2_xor3v1x2_0_bn totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1234 totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_1_diff2_2_xor3v1x2_0_bn totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1235 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_in_a totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1236 totdiff3_1_diff2_2_xor3v1x2_0_bn totdiff3_1_diff2_2_in_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1237 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_xor3v1x2_0_bn totdiff3_0_mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1238 totdiff3_1_diff2_2_xor3v1x2_0_a_11_12# totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1239 totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_xor3v1x2_0_a_11_12# totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1240 totdiff3_1_diff2_2_xor3v1x2_0_a_28_12# totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_mux_0_a2 totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1241 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_diff2_2_xor3v1x2_0_a_28_12# totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1242 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1243 totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_in_c totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1244 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_in_c totdiff3_1_mux_0_a2 totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1245 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1246 totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_diff2_2_in_c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1247 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_in_c totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1248 totdiff3_1_diff2_2_xor3v1x2_0_a_115_7# totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1249 totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_1_diff2_2_xor3v1x2_0_bn totdiff3_1_diff2_2_xor3v1x2_0_a_115_7# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1250 totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1251 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_in_a totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1252 totdiff3_1_diff2_2_xor3v1x2_0_bn totdiff3_1_diff2_2_in_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1253 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_an2v0x2_2_zn totdiff3_1_diff2_2_in_2c totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1254 totdiff3_1_diff2_1_an2v0x2_2_zn totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1255 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_in_2c totdiff3_1_diff2_1_an2v0x2_2_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1256 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_an2v0x2_2_zn totdiff3_1_diff2_2_in_2c totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1257 totdiff3_1_diff2_1_an2v0x2_2_a_24_13# totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1258 totdiff3_1_diff2_1_an2v0x2_2_zn totdiff3_1_diff2_1_in_2c totdiff3_1_diff2_1_an2v0x2_2_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1259 totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_mux_0_b1 totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1260 totdiff3_1_mux_0_b1 totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1261 totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_1_mux_0_b1 totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1262 totdiff3_1_mux_0_b1 totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1263 totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_diff2_1_in_2c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1264 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_in_2c totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1265 totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1266 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1267 totdiff3_1_diff2_1_xor2v2x2_0_a_13_13# totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1268 totdiff3_1_mux_0_b1 totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_diff2_1_xor2v2x2_0_a_13_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1269 totdiff3_1_diff2_1_xor2v2x2_0_a_30_13# totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_mux_0_b1 totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1270 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_1_diff2_1_xor2v2x2_0_a_30_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1271 totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_diff2_1_in_2c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1272 totdiff3_1_mux_0_b1 totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1273 totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_1_diff2_1_in_2c totdiff3_1_mux_0_b1 totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1274 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1275 totdiff3_1_diff2_2_in_c totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1276 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_1_diff2_2_in_c totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1277 totdiff3_1_diff2_1_or2v0x3_0_a_31_39# totdiff3_1_diff2_1_an2v0x2_1_z totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1278 totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_1_diff2_1_an2v0x2_0_z totdiff3_1_diff2_1_or2v0x3_0_a_31_39# totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1279 totdiff3_1_diff2_1_or2v0x3_0_a_48_39# totdiff3_1_diff2_1_an2v0x2_0_z totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1280 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_an2v0x2_1_z totdiff3_1_diff2_1_or2v0x3_0_a_48_39# totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1281 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_1_diff2_2_in_c totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1282 totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_1_diff2_1_an2v0x2_1_z totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1283 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_an2v0x2_0_z totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1284 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_an2v0x2_1_zn totdiff3_1_diff2_1_an2v0x2_1_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1285 totdiff3_1_diff2_1_an2v0x2_1_zn totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1286 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_an2v0x2_1_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1287 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_an2v0x2_1_zn totdiff3_1_diff2_1_an2v0x2_1_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1288 totdiff3_1_diff2_1_an2v0x2_1_a_24_13# totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1289 totdiff3_1_diff2_1_an2v0x2_1_zn totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_an2v0x2_1_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1290 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_an2v0x2_0_zn totdiff3_1_diff2_1_an2v0x2_0_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1291 totdiff3_1_diff2_1_an2v0x2_0_zn totdiff3_1_diff2_1_in_c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1292 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_an2v0x2_0_b totdiff3_1_diff2_1_an2v0x2_0_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1293 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_an2v0x2_0_zn totdiff3_1_diff2_1_an2v0x2_0_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1294 totdiff3_1_diff2_1_an2v0x2_0_a_24_13# totdiff3_1_diff2_1_in_c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1295 totdiff3_1_diff2_1_an2v0x2_0_zn totdiff3_1_diff2_1_an2v0x2_0_b totdiff3_1_diff2_1_an2v0x2_0_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1296 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_xnr2v8x05_0_zn totdiff3_1_diff2_1_an2v0x2_0_b totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1297 totdiff3_1_diff2_1_xnr2v8x05_0_an totdiff3_1_diff2_1_in_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1298 totdiff3_1_diff2_1_xnr2v8x05_0_zn totdiff3_1_diff2_1_xnr2v8x05_0_bn totdiff3_1_diff2_1_xnr2v8x05_0_an totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1299 totdiff3_1_diff2_1_xnr2v8x05_0_ai totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_xnr2v8x05_0_zn totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1300 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_xnr2v8x05_0_an totdiff3_1_diff2_1_xnr2v8x05_0_ai totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1301 totdiff3_1_diff2_1_xnr2v8x05_0_bn totdiff3_1_diff2_1_in_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1302 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xnr2v8x05_0_zn totdiff3_1_diff2_1_an2v0x2_0_b totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1303 totdiff3_1_diff2_1_xnr2v8x05_0_an totdiff3_1_diff2_1_in_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1304 totdiff3_1_diff2_1_xnr2v8x05_0_zn totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_xnr2v8x05_0_an totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1305 totdiff3_1_diff2_1_xnr2v8x05_0_ai totdiff3_1_diff2_1_xnr2v8x05_0_bn totdiff3_1_diff2_1_xnr2v8x05_0_zn totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1306 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xnr2v8x05_0_an totdiff3_1_diff2_1_xnr2v8x05_0_ai totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1307 totdiff3_1_diff2_1_xnr2v8x05_0_bn totdiff3_1_diff2_1_in_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1308 totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_1_mux_0_a1 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1309 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1310 totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_1_mux_0_a1 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1311 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1312 totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_mux_0_a1 totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1313 totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1314 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_mux_0_a1 totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1315 totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1316 totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_diff2_1_in_c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1317 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_in_c totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_0_mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1318 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1319 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1320 totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1321 totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1322 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_in_a totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1323 totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_1_diff2_1_in_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1324 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_0_mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1325 totdiff3_1_diff2_1_xor3v1x2_0_a_11_12# totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1326 totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_xor3v1x2_0_a_11_12# totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1327 totdiff3_1_diff2_1_xor3v1x2_0_a_28_12# totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_mux_0_a1 totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1328 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_diff2_1_xor3v1x2_0_a_28_12# totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1329 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1330 totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_in_c totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1331 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_in_c totdiff3_1_mux_0_a1 totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1332 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1333 totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_diff2_1_in_c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1334 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_in_c totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1335 totdiff3_1_diff2_1_xor3v1x2_0_a_115_7# totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1336 totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_1_diff2_1_xor3v1x2_0_a_115_7# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1337 totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1338 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_in_a totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1339 totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_1_diff2_1_in_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1340 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_an2v0x2_2_zn totdiff3_1_diff2_1_in_2c totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1341 totdiff3_1_diff2_0_an2v0x2_2_zn totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1342 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_an2v0x2_2_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1343 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_an2v0x2_2_zn totdiff3_1_diff2_1_in_2c totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1344 totdiff3_1_diff2_0_an2v0x2_2_a_24_13# totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1345 totdiff3_1_diff2_0_an2v0x2_2_zn totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_an2v0x2_2_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1346 totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_1_mux_0_b0 totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1347 totdiff3_1_mux_0_b0 totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1348 totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_1_mux_0_b0 totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1349 totdiff3_1_mux_0_b0 totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1350 totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1351 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1352 totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1353 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1354 totdiff3_1_diff2_0_xor2v2x2_0_a_13_13# totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1355 totdiff3_1_mux_0_b0 totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_1_diff2_0_xor2v2x2_0_a_13_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1356 totdiff3_1_diff2_0_xor2v2x2_0_a_30_13# totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_1_mux_0_b0 totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1357 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_1_diff2_0_xor2v2x2_0_a_30_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1358 totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_vdd totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1359 totdiff3_1_mux_0_b0 totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1360 totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_0_mux_0_vdd totdiff3_1_mux_0_b0 totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1361 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1362 totdiff3_1_diff2_1_in_c totdiff3_1_diff2_0_or2v0x3_0_zn totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1363 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_or2v0x3_0_zn totdiff3_1_diff2_1_in_c totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1364 totdiff3_1_diff2_0_or2v0x3_0_a_31_39# totdiff3_1_diff2_0_an2v0x2_1_z totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1365 totdiff3_1_diff2_0_or2v0x3_0_zn totdiff3_1_diff2_0_an2v0x2_0_z totdiff3_1_diff2_0_or2v0x3_0_a_31_39# totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1366 totdiff3_1_diff2_0_or2v0x3_0_a_48_39# totdiff3_1_diff2_0_an2v0x2_0_z totdiff3_1_diff2_0_or2v0x3_0_zn totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1367 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_an2v0x2_1_z totdiff3_1_diff2_0_or2v0x3_0_a_48_39# totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1368 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_or2v0x3_0_zn totdiff3_1_diff2_1_in_c totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1369 totdiff3_1_diff2_0_or2v0x3_0_zn totdiff3_1_diff2_0_an2v0x2_1_z totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1370 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_an2v0x2_0_z totdiff3_1_diff2_0_or2v0x3_0_zn totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1371 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_an2v0x2_1_zn totdiff3_1_diff2_0_an2v0x2_1_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1372 totdiff3_1_diff2_0_an2v0x2_1_zn totdiff3_1_diff2_0_an2v0x2_1_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1373 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_an2v0x2_1_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1374 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_an2v0x2_1_zn totdiff3_1_diff2_0_an2v0x2_1_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1375 totdiff3_1_diff2_0_an2v0x2_1_a_24_13# totdiff3_1_diff2_0_an2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1376 totdiff3_1_diff2_0_an2v0x2_1_zn totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_an2v0x2_1_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1377 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_an2v0x2_0_zn totdiff3_1_diff2_0_an2v0x2_0_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1378 totdiff3_1_diff2_0_an2v0x2_0_zn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1379 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_an2v0x2_0_b totdiff3_1_diff2_0_an2v0x2_0_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1380 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_an2v0x2_0_zn totdiff3_1_diff2_0_an2v0x2_0_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1381 totdiff3_1_diff2_0_an2v0x2_0_a_24_13# totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1382 totdiff3_1_diff2_0_an2v0x2_0_zn totdiff3_1_diff2_0_an2v0x2_0_b totdiff3_1_diff2_0_an2v0x2_0_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1383 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_xnr2v8x05_0_zn totdiff3_1_diff2_0_an2v0x2_0_b totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1384 totdiff3_1_diff2_0_xnr2v8x05_0_an totdiff3_1_diff2_0_in_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1385 totdiff3_1_diff2_0_xnr2v8x05_0_zn totdiff3_1_diff2_0_xnr2v8x05_0_bn totdiff3_1_diff2_0_xnr2v8x05_0_an totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1386 totdiff3_1_diff2_0_xnr2v8x05_0_ai totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_xnr2v8x05_0_zn totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1387 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_xnr2v8x05_0_an totdiff3_1_diff2_0_xnr2v8x05_0_ai totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1388 totdiff3_1_diff2_0_xnr2v8x05_0_bn totdiff3_1_diff2_0_in_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1389 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xnr2v8x05_0_zn totdiff3_1_diff2_0_an2v0x2_0_b totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1390 totdiff3_1_diff2_0_xnr2v8x05_0_an totdiff3_1_diff2_0_in_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1391 totdiff3_1_diff2_0_xnr2v8x05_0_zn totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_xnr2v8x05_0_an totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1392 totdiff3_1_diff2_0_xnr2v8x05_0_ai totdiff3_1_diff2_0_xnr2v8x05_0_bn totdiff3_1_diff2_0_xnr2v8x05_0_zn totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1393 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xnr2v8x05_0_an totdiff3_1_diff2_0_xnr2v8x05_0_ai totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1394 totdiff3_1_diff2_0_xnr2v8x05_0_bn totdiff3_1_diff2_0_in_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1395 totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_1_mux_0_a0 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1396 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1397 totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_1_mux_0_a0 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1398 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1399 totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_mux_0_a0 totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1400 totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1401 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_1_mux_0_a0 totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1402 totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1403 totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1404 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1405 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1406 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1407 totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_1_diff2_0_an2v0x2_1_a totdiff3_1_diff2_0_xor3v1x2_0_bn totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1408 totdiff3_1_diff2_0_an2v0x2_1_a totdiff3_1_diff2_0_xor3v1x2_0_bn totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1409 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_in_a totdiff3_1_diff2_0_an2v0x2_1_a totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1410 totdiff3_1_diff2_0_xor3v1x2_0_bn totdiff3_1_diff2_0_in_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1411 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_xor3v1x2_0_bn totdiff3_0_mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1412 totdiff3_1_diff2_0_xor3v1x2_0_a_11_12# totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1413 totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_diff2_0_xor3v1x2_0_a_11_12# totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1414 totdiff3_1_diff2_0_xor3v1x2_0_a_28_12# totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_mux_0_a0 totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1415 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_1_diff2_0_xor3v1x2_0_a_28_12# totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1416 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1417 totdiff3_1_mux_0_a0 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1418 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_gnd totdiff3_1_mux_0_a0 totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1419 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1420 totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1421 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1422 totdiff3_1_diff2_0_xor3v1x2_0_a_115_7# totdiff3_1_diff2_0_an2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1423 totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_1_diff2_0_xor3v1x2_0_bn totdiff3_1_diff2_0_xor3v1x2_0_a_115_7# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1424 totdiff3_1_diff2_0_an2v0x2_1_a totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1425 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_in_a totdiff3_1_diff2_0_an2v0x2_1_a totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1426 totdiff3_1_diff2_0_xor3v1x2_0_bn totdiff3_1_diff2_0_in_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1427 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_2_zn comp_0_an3v0x2_2_c totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1428 totdiff3_0_mux_0_mxn2v0x1_2_a_21_50# totdiff3_0_mux_0_a2 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1429 totdiff3_0_mux_0_mxn2v0x1_2_zn totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_2_a_21_50# totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1430 totdiff3_0_mux_0_mxn2v0x1_2_a_38_50# totdiff3_0_mux_0_mxn2v0x1_2_sn totdiff3_0_mux_0_mxn2v0x1_2_zn totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1431 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_b2 totdiff3_0_mux_0_mxn2v0x1_2_a_38_50# totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1432 totdiff3_0_mux_0_mxn2v0x1_2_sn totdiff3_0_mux_0_s totdiff3_0_mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1433 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_2_zn comp_0_an3v0x2_2_c totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1434 totdiff3_0_mux_0_mxn2v0x1_2_a_21_12# totdiff3_0_mux_0_a2 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1435 totdiff3_0_mux_0_mxn2v0x1_2_zn totdiff3_0_mux_0_mxn2v0x1_2_sn totdiff3_0_mux_0_mxn2v0x1_2_a_21_12# totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1436 totdiff3_0_mux_0_mxn2v0x1_2_a_38_12# totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_2_zn totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1437 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_b2 totdiff3_0_mux_0_mxn2v0x1_2_a_38_12# totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1438 totdiff3_0_mux_0_mxn2v0x1_2_sn totdiff3_0_mux_0_s totdiff3_0_mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1439 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_1_zn comp_0_an3v0x2_0_b totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1440 totdiff3_0_mux_0_mxn2v0x1_1_a_21_50# totdiff3_0_mux_0_a1 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1441 totdiff3_0_mux_0_mxn2v0x1_1_zn totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_1_a_21_50# totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1442 totdiff3_0_mux_0_mxn2v0x1_1_a_38_50# totdiff3_0_mux_0_mxn2v0x1_1_sn totdiff3_0_mux_0_mxn2v0x1_1_zn totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1443 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_b1 totdiff3_0_mux_0_mxn2v0x1_1_a_38_50# totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1444 totdiff3_0_mux_0_mxn2v0x1_1_sn totdiff3_0_mux_0_s totdiff3_0_mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1445 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_1_zn comp_0_an3v0x2_0_b totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1446 totdiff3_0_mux_0_mxn2v0x1_1_a_21_12# totdiff3_0_mux_0_a1 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1447 totdiff3_0_mux_0_mxn2v0x1_1_zn totdiff3_0_mux_0_mxn2v0x1_1_sn totdiff3_0_mux_0_mxn2v0x1_1_a_21_12# totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1448 totdiff3_0_mux_0_mxn2v0x1_1_a_38_12# totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_1_zn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1449 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_b1 totdiff3_0_mux_0_mxn2v0x1_1_a_38_12# totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1450 totdiff3_0_mux_0_mxn2v0x1_1_sn totdiff3_0_mux_0_s totdiff3_0_mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1451 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_0_zn comp_0_an3v0x2_2_a totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1452 totdiff3_0_mux_0_mxn2v0x1_0_a_21_50# totdiff3_0_mux_0_a0 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1453 totdiff3_0_mux_0_mxn2v0x1_0_zn totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_0_a_21_50# totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1454 totdiff3_0_mux_0_mxn2v0x1_0_a_38_50# totdiff3_0_mux_0_mxn2v0x1_0_sn totdiff3_0_mux_0_mxn2v0x1_0_zn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1455 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_b0 totdiff3_0_mux_0_mxn2v0x1_0_a_38_50# totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1456 totdiff3_0_mux_0_mxn2v0x1_0_sn totdiff3_0_mux_0_s totdiff3_0_mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1457 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_0_zn comp_0_an3v0x2_2_a totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1458 totdiff3_0_mux_0_mxn2v0x1_0_a_21_12# totdiff3_0_mux_0_a0 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1459 totdiff3_0_mux_0_mxn2v0x1_0_zn totdiff3_0_mux_0_mxn2v0x1_0_sn totdiff3_0_mux_0_mxn2v0x1_0_a_21_12# totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1460 totdiff3_0_mux_0_mxn2v0x1_0_a_38_12# totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_0_zn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1461 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_b0 totdiff3_0_mux_0_mxn2v0x1_0_a_38_12# totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1462 totdiff3_0_mux_0_mxn2v0x1_0_sn totdiff3_0_mux_0_s totdiff3_0_mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1463 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_an2v0x2_2_zn totdiff3_0_diff2_2_an2v0x2_2_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1464 totdiff3_0_diff2_2_an2v0x2_2_zn totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1465 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_in_2c totdiff3_0_diff2_2_an2v0x2_2_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1466 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_2_zn totdiff3_0_diff2_2_an2v0x2_2_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1467 totdiff3_0_diff2_2_an2v0x2_2_a_24_13# totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1468 totdiff3_0_diff2_2_an2v0x2_2_zn totdiff3_0_diff2_2_in_2c totdiff3_0_diff2_2_an2v0x2_2_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1469 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_mux_0_b2 totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1470 totdiff3_0_mux_0_b2 totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1471 totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_b2 totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1472 totdiff3_0_mux_0_b2 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1473 totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_diff2_2_in_2c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1474 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_in_2c totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1475 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1476 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1477 totdiff3_0_diff2_2_xor2v2x2_0_a_13_13# totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1478 totdiff3_0_mux_0_b2 totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_diff2_2_xor2v2x2_0_a_13_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1479 totdiff3_0_diff2_2_xor2v2x2_0_a_30_13# totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_mux_0_b2 totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1480 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_diff2_2_xor2v2x2_0_a_30_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1481 totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_diff2_2_in_2c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1482 totdiff3_0_mux_0_b2 totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1483 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_diff2_2_in_2c totdiff3_0_mux_0_b2 totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1484 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1485 totdiff3_0_mux_0_s totdiff3_0_diff2_2_or2v0x3_0_zn totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1486 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_or2v0x3_0_zn totdiff3_0_mux_0_s totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1487 totdiff3_0_diff2_2_or2v0x3_0_a_31_39# totdiff3_0_diff2_2_an2v0x2_1_z totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1488 totdiff3_0_diff2_2_or2v0x3_0_zn totdiff3_0_diff2_2_an2v0x2_0_z totdiff3_0_diff2_2_or2v0x3_0_a_31_39# totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1489 totdiff3_0_diff2_2_or2v0x3_0_a_48_39# totdiff3_0_diff2_2_an2v0x2_0_z totdiff3_0_diff2_2_or2v0x3_0_zn totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1490 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_an2v0x2_1_z totdiff3_0_diff2_2_or2v0x3_0_a_48_39# totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1491 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_or2v0x3_0_zn totdiff3_0_mux_0_s totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1492 totdiff3_0_diff2_2_or2v0x3_0_zn totdiff3_0_diff2_2_an2v0x2_1_z totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1493 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_0_z totdiff3_0_diff2_2_or2v0x3_0_zn totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1494 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_an2v0x2_1_zn totdiff3_0_diff2_2_an2v0x2_1_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1495 totdiff3_0_diff2_2_an2v0x2_1_zn totdiff3_0_diff2_2_an2v0x2_1_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1496 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_an2v0x2_1_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1497 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_1_zn totdiff3_0_diff2_2_an2v0x2_1_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1498 totdiff3_0_diff2_2_an2v0x2_1_a_24_13# totdiff3_0_diff2_2_an2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1499 totdiff3_0_diff2_2_an2v0x2_1_zn totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_an2v0x2_1_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1500 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_an2v0x2_0_zn totdiff3_0_diff2_2_an2v0x2_0_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1501 totdiff3_0_diff2_2_an2v0x2_0_zn totdiff3_0_diff2_2_in_c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1502 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_an2v0x2_0_b totdiff3_0_diff2_2_an2v0x2_0_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1503 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_0_zn totdiff3_0_diff2_2_an2v0x2_0_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1504 totdiff3_0_diff2_2_an2v0x2_0_a_24_13# totdiff3_0_diff2_2_in_c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1505 totdiff3_0_diff2_2_an2v0x2_0_zn totdiff3_0_diff2_2_an2v0x2_0_b totdiff3_0_diff2_2_an2v0x2_0_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1506 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_xnr2v8x05_0_zn totdiff3_0_diff2_2_an2v0x2_0_b totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1507 totdiff3_0_diff2_2_xnr2v8x05_0_an totdiff3_0_diff2_2_in_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1508 totdiff3_0_diff2_2_xnr2v8x05_0_zn totdiff3_0_diff2_2_xnr2v8x05_0_bn totdiff3_0_diff2_2_xnr2v8x05_0_an totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1509 totdiff3_0_diff2_2_xnr2v8x05_0_ai totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_xnr2v8x05_0_zn totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1510 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_xnr2v8x05_0_an totdiff3_0_diff2_2_xnr2v8x05_0_ai totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1511 totdiff3_0_diff2_2_xnr2v8x05_0_bn totdiff3_0_diff2_2_in_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1512 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xnr2v8x05_0_zn totdiff3_0_diff2_2_an2v0x2_0_b totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1513 totdiff3_0_diff2_2_xnr2v8x05_0_an totdiff3_0_diff2_2_in_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1514 totdiff3_0_diff2_2_xnr2v8x05_0_zn totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_xnr2v8x05_0_an totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1515 totdiff3_0_diff2_2_xnr2v8x05_0_ai totdiff3_0_diff2_2_xnr2v8x05_0_bn totdiff3_0_diff2_2_xnr2v8x05_0_zn totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1516 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xnr2v8x05_0_an totdiff3_0_diff2_2_xnr2v8x05_0_ai totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1517 totdiff3_0_diff2_2_xnr2v8x05_0_bn totdiff3_0_diff2_2_in_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1518 totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_a2 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1519 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1520 totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_a2 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1521 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1522 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_a2 totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1523 totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1524 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_mux_0_a2 totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1525 totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1526 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_in_c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1527 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_in_c totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1528 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1529 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1530 totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_diff2_2_an2v0x2_1_a totdiff3_0_diff2_2_xor3v1x2_0_bn totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1531 totdiff3_0_diff2_2_an2v0x2_1_a totdiff3_0_diff2_2_xor3v1x2_0_bn totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1532 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_in_a totdiff3_0_diff2_2_an2v0x2_1_a totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1533 totdiff3_0_diff2_2_xor3v1x2_0_bn totdiff3_0_diff2_2_in_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1534 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_xor3v1x2_0_bn totdiff3_0_mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1535 totdiff3_0_diff2_2_xor3v1x2_0_a_11_12# totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1536 totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_xor3v1x2_0_a_11_12# totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1537 totdiff3_0_diff2_2_xor3v1x2_0_a_28_12# totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_a2 totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1538 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_xor3v1x2_0_a_28_12# totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1539 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1540 totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_in_c totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1541 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_in_c totdiff3_0_mux_0_a2 totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1542 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1543 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_in_c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1544 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_in_c totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1545 totdiff3_0_diff2_2_xor3v1x2_0_a_115_7# totdiff3_0_diff2_2_an2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1546 totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_diff2_2_xor3v1x2_0_bn totdiff3_0_diff2_2_xor3v1x2_0_a_115_7# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1547 totdiff3_0_diff2_2_an2v0x2_1_a totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1548 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_in_a totdiff3_0_diff2_2_an2v0x2_1_a totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1549 totdiff3_0_diff2_2_xor3v1x2_0_bn totdiff3_0_diff2_2_in_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1550 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_2_zn totdiff3_0_diff2_2_in_2c totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1551 totdiff3_0_diff2_1_an2v0x2_2_zn totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1552 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_in_2c totdiff3_0_diff2_1_an2v0x2_2_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1553 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_2_zn totdiff3_0_diff2_2_in_2c totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1554 totdiff3_0_diff2_1_an2v0x2_2_a_24_13# totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1555 totdiff3_0_diff2_1_an2v0x2_2_zn totdiff3_0_diff2_1_in_2c totdiff3_0_diff2_1_an2v0x2_2_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1556 totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_mux_0_b1 totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1557 totdiff3_0_mux_0_b1 totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1558 totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_mux_0_b1 totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1559 totdiff3_0_mux_0_b1 totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1560 totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_diff2_1_in_2c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1561 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_in_2c totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1562 totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1563 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1564 totdiff3_0_diff2_1_xor2v2x2_0_a_13_13# totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1565 totdiff3_0_mux_0_b1 totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_diff2_1_xor2v2x2_0_a_13_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1566 totdiff3_0_diff2_1_xor2v2x2_0_a_30_13# totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_mux_0_b1 totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1567 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_diff2_1_xor2v2x2_0_a_30_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1568 totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_diff2_1_in_2c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1569 totdiff3_0_mux_0_b1 totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1570 totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_diff2_1_in_2c totdiff3_0_mux_0_b1 totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1571 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1572 totdiff3_0_diff2_2_in_c totdiff3_0_diff2_1_or2v0x3_0_zn totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1573 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_or2v0x3_0_zn totdiff3_0_diff2_2_in_c totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1574 totdiff3_0_diff2_1_or2v0x3_0_a_31_39# totdiff3_0_diff2_1_an2v0x2_1_z totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1575 totdiff3_0_diff2_1_or2v0x3_0_zn totdiff3_0_diff2_1_an2v0x2_0_z totdiff3_0_diff2_1_or2v0x3_0_a_31_39# totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1576 totdiff3_0_diff2_1_or2v0x3_0_a_48_39# totdiff3_0_diff2_1_an2v0x2_0_z totdiff3_0_diff2_1_or2v0x3_0_zn totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1577 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_1_z totdiff3_0_diff2_1_or2v0x3_0_a_48_39# totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1578 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_or2v0x3_0_zn totdiff3_0_diff2_2_in_c totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1579 totdiff3_0_diff2_1_or2v0x3_0_zn totdiff3_0_diff2_1_an2v0x2_1_z totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1580 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_0_z totdiff3_0_diff2_1_or2v0x3_0_zn totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1581 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_1_zn totdiff3_0_diff2_1_an2v0x2_1_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1582 totdiff3_0_diff2_1_an2v0x2_1_zn totdiff3_0_diff2_1_an2v0x2_1_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1583 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_an2v0x2_1_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1584 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_1_zn totdiff3_0_diff2_1_an2v0x2_1_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1585 totdiff3_0_diff2_1_an2v0x2_1_a_24_13# totdiff3_0_diff2_1_an2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1586 totdiff3_0_diff2_1_an2v0x2_1_zn totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_an2v0x2_1_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1587 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_0_zn totdiff3_0_diff2_1_an2v0x2_0_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1588 totdiff3_0_diff2_1_an2v0x2_0_zn totdiff3_0_diff2_1_in_c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1589 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_0_b totdiff3_0_diff2_1_an2v0x2_0_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1590 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_0_zn totdiff3_0_diff2_1_an2v0x2_0_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1591 totdiff3_0_diff2_1_an2v0x2_0_a_24_13# totdiff3_0_diff2_1_in_c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1592 totdiff3_0_diff2_1_an2v0x2_0_zn totdiff3_0_diff2_1_an2v0x2_0_b totdiff3_0_diff2_1_an2v0x2_0_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1593 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_xnr2v8x05_0_zn totdiff3_0_diff2_1_an2v0x2_0_b totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1594 totdiff3_0_diff2_1_xnr2v8x05_0_an totdiff3_0_diff2_1_in_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1595 totdiff3_0_diff2_1_xnr2v8x05_0_zn totdiff3_0_diff2_1_xnr2v8x05_0_bn totdiff3_0_diff2_1_xnr2v8x05_0_an totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1596 totdiff3_0_diff2_1_xnr2v8x05_0_ai totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_xnr2v8x05_0_zn totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1597 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_xnr2v8x05_0_an totdiff3_0_diff2_1_xnr2v8x05_0_ai totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1598 totdiff3_0_diff2_1_xnr2v8x05_0_bn totdiff3_0_diff2_1_in_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1599 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xnr2v8x05_0_zn totdiff3_0_diff2_1_an2v0x2_0_b totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1600 totdiff3_0_diff2_1_xnr2v8x05_0_an totdiff3_0_diff2_1_in_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1601 totdiff3_0_diff2_1_xnr2v8x05_0_zn totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_xnr2v8x05_0_an totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1602 totdiff3_0_diff2_1_xnr2v8x05_0_ai totdiff3_0_diff2_1_xnr2v8x05_0_bn totdiff3_0_diff2_1_xnr2v8x05_0_zn totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1603 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xnr2v8x05_0_an totdiff3_0_diff2_1_xnr2v8x05_0_ai totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1604 totdiff3_0_diff2_1_xnr2v8x05_0_bn totdiff3_0_diff2_1_in_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1605 totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_a1 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1606 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1607 totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_a1 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1608 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1609 totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_a1 totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1610 totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1611 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_mux_0_a1 totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1612 totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1613 totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_diff2_1_in_c totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1614 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_in_c totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1615 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1616 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1617 totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_diff2_1_an2v0x2_1_a totdiff3_0_diff2_1_xor3v1x2_0_bn totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1618 totdiff3_0_diff2_1_an2v0x2_1_a totdiff3_0_diff2_1_xor3v1x2_0_bn totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1619 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_in_a totdiff3_0_diff2_1_an2v0x2_1_a totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1620 totdiff3_0_diff2_1_xor3v1x2_0_bn totdiff3_0_diff2_1_in_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1621 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_xor3v1x2_0_bn totdiff3_0_mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1622 totdiff3_0_diff2_1_xor3v1x2_0_a_11_12# totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1623 totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_xor3v1x2_0_a_11_12# totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1624 totdiff3_0_diff2_1_xor3v1x2_0_a_28_12# totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_a1 totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1625 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_diff2_1_xor3v1x2_0_a_28_12# totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1626 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1627 totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_in_c totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1628 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_in_c totdiff3_0_mux_0_a1 totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1629 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1630 totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_diff2_1_in_c totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1631 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_in_c totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1632 totdiff3_0_diff2_1_xor3v1x2_0_a_115_7# totdiff3_0_diff2_1_an2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1633 totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_diff2_1_xor3v1x2_0_bn totdiff3_0_diff2_1_xor3v1x2_0_a_115_7# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1634 totdiff3_0_diff2_1_an2v0x2_1_a totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1635 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_in_a totdiff3_0_diff2_1_an2v0x2_1_a totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1636 totdiff3_0_diff2_1_xor3v1x2_0_bn totdiff3_0_diff2_1_in_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1637 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_2_zn totdiff3_0_diff2_1_in_2c totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1638 totdiff3_0_diff2_0_an2v0x2_2_zn totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1639 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_2_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1640 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_2_zn totdiff3_0_diff2_1_in_2c totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1641 totdiff3_0_diff2_0_an2v0x2_2_a_24_13# totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1642 totdiff3_0_diff2_0_an2v0x2_2_zn totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_2_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1643 totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_b0 totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1644 totdiff3_0_mux_0_b0 totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1645 totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_mux_0_b0 totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1646 totdiff3_0_mux_0_b0 totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1647 totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1648 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1649 totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1650 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1651 totdiff3_0_diff2_0_xor2v2x2_0_a_13_13# totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1652 totdiff3_0_mux_0_b0 totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_diff2_0_xor2v2x2_0_a_13_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1653 totdiff3_0_diff2_0_xor2v2x2_0_a_30_13# totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_b0 totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1654 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_diff2_0_xor2v2x2_0_a_30_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1655 totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_vdd totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1656 totdiff3_0_mux_0_b0 totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1657 totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_mux_0_vdd totdiff3_0_mux_0_b0 totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1658 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1659 totdiff3_0_diff2_1_in_c totdiff3_0_diff2_0_or2v0x3_0_zn totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1660 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_or2v0x3_0_zn totdiff3_0_diff2_1_in_c totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1661 totdiff3_0_diff2_0_or2v0x3_0_a_31_39# totdiff3_0_diff2_0_an2v0x2_1_z totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1662 totdiff3_0_diff2_0_or2v0x3_0_zn totdiff3_0_diff2_0_an2v0x2_0_z totdiff3_0_diff2_0_or2v0x3_0_a_31_39# totdiff3_0_mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1663 totdiff3_0_diff2_0_or2v0x3_0_a_48_39# totdiff3_0_diff2_0_an2v0x2_0_z totdiff3_0_diff2_0_or2v0x3_0_zn totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1664 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_1_z totdiff3_0_diff2_0_or2v0x3_0_a_48_39# totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1665 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_or2v0x3_0_zn totdiff3_0_diff2_1_in_c totdiff3_0_mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1666 totdiff3_0_diff2_0_or2v0x3_0_zn totdiff3_0_diff2_0_an2v0x2_1_z totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1667 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_0_z totdiff3_0_diff2_0_or2v0x3_0_zn totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1668 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_1_zn totdiff3_0_diff2_0_an2v0x2_1_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1669 totdiff3_0_diff2_0_an2v0x2_1_zn totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1670 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_an2v0x2_1_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1671 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_1_zn totdiff3_0_diff2_0_an2v0x2_1_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1672 totdiff3_0_diff2_0_an2v0x2_1_a_24_13# totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1673 totdiff3_0_diff2_0_an2v0x2_1_zn totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_an2v0x2_1_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1674 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_0_zn totdiff3_0_diff2_0_an2v0x2_0_z totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1675 totdiff3_0_diff2_0_an2v0x2_0_zn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1676 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_0_b totdiff3_0_diff2_0_an2v0x2_0_zn totdiff3_0_mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1677 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_0_zn totdiff3_0_diff2_0_an2v0x2_0_z totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1678 totdiff3_0_diff2_0_an2v0x2_0_a_24_13# totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1679 totdiff3_0_diff2_0_an2v0x2_0_zn totdiff3_0_diff2_0_an2v0x2_0_b totdiff3_0_diff2_0_an2v0x2_0_a_24_13# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1680 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xnr2v8x05_0_zn totdiff3_0_diff2_0_an2v0x2_0_b totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1681 totdiff3_0_diff2_0_xnr2v8x05_0_an totdiff3_0_diff2_0_in_a totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1682 totdiff3_0_diff2_0_xnr2v8x05_0_zn totdiff3_0_diff2_0_xnr2v8x05_0_bn totdiff3_0_diff2_0_xnr2v8x05_0_an totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1683 totdiff3_0_diff2_0_xnr2v8x05_0_ai totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_xnr2v8x05_0_zn totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1684 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xnr2v8x05_0_an totdiff3_0_diff2_0_xnr2v8x05_0_ai totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1685 totdiff3_0_diff2_0_xnr2v8x05_0_bn totdiff3_0_diff2_0_in_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1686 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xnr2v8x05_0_zn totdiff3_0_diff2_0_an2v0x2_0_b totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1687 totdiff3_0_diff2_0_xnr2v8x05_0_an totdiff3_0_diff2_0_in_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1688 totdiff3_0_diff2_0_xnr2v8x05_0_zn totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_xnr2v8x05_0_an totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1689 totdiff3_0_diff2_0_xnr2v8x05_0_ai totdiff3_0_diff2_0_xnr2v8x05_0_bn totdiff3_0_diff2_0_xnr2v8x05_0_zn totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1690 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xnr2v8x05_0_an totdiff3_0_diff2_0_xnr2v8x05_0_ai totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1691 totdiff3_0_diff2_0_xnr2v8x05_0_bn totdiff3_0_diff2_0_in_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1692 totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_a0 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1693 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1694 totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_a0 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1695 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1696 totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_a0 totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1697 totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1698 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_a0 totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1699 totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1700 totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1701 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1702 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1703 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1704 totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1705 totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1706 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_in_a totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1707 totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_diff2_0_in_b totdiff3_0_mux_0_vdd totdiff3_0_mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1708 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1709 totdiff3_0_diff2_0_xor3v1x2_0_a_11_12# totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1710 totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_diff2_0_xor3v1x2_0_a_11_12# totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1711 totdiff3_0_diff2_0_xor3v1x2_0_a_28_12# totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_a0 totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1712 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_diff2_0_xor3v1x2_0_a_28_12# totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1713 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1714 totdiff3_0_mux_0_a0 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1715 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_a0 totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1716 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1717 totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1718 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1719 totdiff3_0_diff2_0_xor3v1x2_0_a_115_7# totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1720 totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_diff2_0_xor3v1x2_0_a_115_7# totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1721 totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1722 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_in_a totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1723 totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_diff2_0_in_b totdiff3_0_mux_0_gnd totdiff3_0_mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
C0 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xor3v1x2_0_bn 15.4fF
C1 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_in_c 34.1fF
C2 totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_xor3v1x2_0_bn 2.6fF
C3 totdiff3_1_diff2_1_in_2c totdiff3_0_mux_0_vdd 34.0fF
C4 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xor2v2x2_0_bn 11.2fF
C5 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_an2v0x2_1_zn 8.9fF
C6 totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_1_diff2_2_in_b 2.0fF
C7 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_2_a 61.1fF
C8 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_0_zn 8.9fF
C9 totdiff3_1_diff2_1_an2v0x2_1_zn totdiff3_0_mux_0_vdd 8.8fF
C10 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_mux_0_a2 4.6fF
C11 totdiff3_1_diff2_2_an2v0x2_1_zn totdiff3_0_mux_0_vdd 8.8fF
C12 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_xor3v1x2_0_bn 9.1fF
C13 comp_0_an2v0x2_1_b totdiff3_0_mux_0_gnd 5.9fF
C14 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_1_z 17.9fF
C15 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_1_mux_0_a2 4.8fF
C16 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_or2v0x3_0_zn 9.0fF
C17 comp_0_an3v0x2_2_c comp_0_nr3v0x2_0_a 2.5fF
C18 totdiff3_1_mux_0_b1 totdiff3_0_mux_0_vdd 13.1fF
C19 comp_0_an2v0x2_3_zn totdiff3_0_mux_0_vdd 8.8fF
C20 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xor3v1x2_0_zn 11.9fF
C21 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xor2v2x2_0_bn 11.2fF
C22 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_an2v0x2_0_z 24.6fF
C23 totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_xor3v1x2_0_cn 4.1fF
C24 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xor2v2x2_0_an 21.6fF
C25 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_in_2c 34.0fF
C26 totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_0_mux_0_gnd 26.1fF
C27 comp_0_iv1v0x4_0_a totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 6.3fF
C28 comp_0_an2v0x2_1_z totdiff3_0_mux_0_vdd 22.0fF
C29 totdiff3_1_diff2_2_or2v0x3_0_zn totdiff3_0_mux_0_vdd 12.7fF
C30 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_xor3v1x2_0_cn 31.6fF
C31 comp_0_an3v0x2_2_a totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 2.3fF
C32 comp_0_an3v0x2_2_a totdiff3_0_mux_0_vdd 42.9fF
C33 totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_xor3v1x2_0_zn 4.6fF
C34 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_a0 14.9fF
C35 comp_0_an3v0x2_2_b comp_0_an2v0x2_0_b 2.5fF
C36 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_in_a 27.8fF
C37 totdiff3_0_diff2_2_in_b totdiff3_0_mux_0_vdd 50.3fF
C38 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_mxn2v0x1_1_zn 9.3fF
C39 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_xor2v2x2_0_an 27.4fF
C40 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_an2v0x2_2_zn 8.9fF
C41 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_gnd 21.6fF
C42 comp_0_an3v0x2_2_c comp_0_an3v0x2_2_w_n4_32# 12.2fF
C43 totdiff3_1_diff2_1_an2v0x2_0_zn totdiff3_0_mux_0_gnd 8.9fF
C44 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_bn 9.1fF
C45 totdiff3_1_diff2_0_xnr2v8x05_0_an totdiff3_0_mux_0_vdd 9.9fF
C46 totdiff3_1_diff2_1_in_2c totdiff3_0_mux_0_gnd 17.5fF
C47 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_xor2v2x2_0_an 25.5fF
C48 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_xor2v2x2_0_bn 17.7fF
C49 totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# 30.3fF
C50 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_an2v0x2_1_z 17.9fF
C51 totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_vdd 59.6fF
C52 comp_0_an2v0x2_1_zn totdiff3_0_mux_0_vdd 8.8fF
C53 comp_0_an3v0x2_1_zn totdiff3_0_mux_0_vdd 4.9fF
C54 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_2_a 25.9fF
C55 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_an2v0x2_1_zn 8.9fF
C56 totdiff3_0_mux_0_mxn2v0x1_1_zn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 8.9fF
C57 comp_0_an3v0x2_2_a totdiff3_1_diff2_1_in_c 9.0fF
C58 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xnr2v8x05_0_zn 4.4fF
C59 totdiff3_1_diff2_2_an2v0x2_1_zn totdiff3_0_mux_0_gnd 8.9fF
C60 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_0_mux_0_vdd 21.4fF
C61 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# comp_0_iv1v0x4_0_a 2.3fF
C62 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_1_z 10.2fF
C63 totdiff3_0_mux_0_b2 totdiff3_0_mux_0_mxn2v0x1_2_zn 2.7fF
C64 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_vdd 25.5fF
C65 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_b1 17.2fF
C66 comp_0_an3v0x2_2_a comp_0_an3v0x2_1_a 6.8fF
C67 totdiff3_0_mux_0_gnd comp_0_an2v0x2_3_zn 8.9fF
C68 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_diff2_0_in_b 4.3fF
C69 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_an2v0x2_0_z 12.8fF
C70 totdiff3_1_diff2_2_xnr2v8x05_0_an totdiff3_0_mux_0_vdd 9.9fF
C71 comp_0_an3v0x2_3_z totdiff3_0_mux_0_vdd 15.4fF
C72 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_in_2c 17.5fF
C73 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# comp_0_iv1v0x4_1_a 2.3fF
C74 totdiff3_0_diff2_2_an2v0x2_2_zn totdiff3_0_mux_0_vdd 8.8fF
C75 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_or2v0x3_0_zn 12.7fF
C76 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_or2v0x3_0_zn 9.0fF
C77 comp_0_an2v0x2_1_z totdiff3_0_mux_0_gnd 8.7fF
C78 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_2_zn 10.3fF
C79 totdiff3_0_diff2_1_in_c totdiff3_0_diff2_1_xnr2v8x05_0_zn 3.1fF
C80 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xor3v1x2_0_cn 18.8fF
C81 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_an2v0x2_0_b 20.5fF
C82 comp_0_an3v0x2_0_b comp_0_an3v0x2_3_zn 3.6fF
C83 comp_0_an3v0x2_2_a totdiff3_0_mux_0_gnd 62.9fF
C84 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_in_b 4.3fF
C85 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_xor3v1x2_0_cn 31.6fF
C86 totdiff3_0_diff2_2_in_b totdiff3_0_mux_0_gnd 60.5fF
C87 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xor2v2x2_0_an 21.6fF
C88 totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_1_diff2_1_in_b 2.6fF
C89 totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_0_mux_0_vdd 12.4fF
C90 comp_0_nr3v0x2_0_a totdiff3_0_mux_0_vdd 4.0fF
C91 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_xor3v1x2_0_cn 31.6fF
C92 totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_0_mux_0_vdd 15.4fF
C93 totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_diff2_1_xor3v1x2_0_cn 2.3fF
C94 totdiff3_1_diff2_0_xnr2v8x05_0_an totdiff3_0_mux_0_gnd 6.8fF
C95 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xor2v2x2_0_an 21.6fF
C96 comp_0_an3v0x2_2_b totdiff3_0_mux_0_vdd 39.7fF
C97 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xor2v2x2_0_bn 11.2fF
C98 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_xor3v1x2_0_bn 15.4fF
C99 comp_0_an3v0x2_3_zn totdiff3_0_mux_0_vdd 10.7fF
C100 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_an2v0x2_2_a 2.3fF
C101 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_an2v0x2_1_z 10.2fF
C102 totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_gnd 25.9fF
C103 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_or2v0x3_0_zn 12.7fF
C104 totdiff3_0_mux_0_gnd comp_0_an2v0x2_1_zn 8.9fF
C105 comp_0_an3v0x2_1_zn totdiff3_0_mux_0_gnd 8.8fF
C106 totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_xor3v1x2_0_zn 4.3fF
C107 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_xor3v1x2_0_zn 18.9fF
C108 comp_0_or3v0x2_0_zn totdiff3_0_mux_0_vdd 9.0fF
C109 totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_xor3v1x2_0_cn 4.1fF
C110 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xnr2v8x05_0_zn 15.0fF
C111 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_0_zn 8.8fF
C112 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_gnd 21.6fF
C113 totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_0_mux_0_a2 4.8fF
C114 totdiff3_1_mux_0_b1 totdiff3_1_mux_0_a1 39.4fF
C115 totdiff3_1_mux_0_s totdiff3_0_mux_0_vdd 7.9fF
C116 comp_0_an3v0x2_2_w_n4_32# totdiff3_0_mux_0_vdd 86.9fF
C117 totdiff3_1_diff2_2_in_a totdiff3_1_diff2_2_an2v0x2_0_zn 2.2fF
C118 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_1_zn 8.8fF
C119 comp_0_an3v0x2_2_b comp_0_an3v0x2_1_a 5.2fF
C120 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_xor3v1x2_0_cn 31.6fF
C121 totdiff3_1_diff2_2_xnr2v8x05_0_an totdiff3_0_mux_0_gnd 5.5fF
C122 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_1_mux_0_mxn2v0x1_0_sn 9.2fF
C123 comp_0_an3v0x2_3_z totdiff3_0_mux_0_gnd 10.6fF
C124 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_in_a 24.6fF
C125 totdiff3_0_mux_0_b2 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# 6.6fF
C126 totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_1_diff2_2_xor3v1x2_0_bn 2.4fF
C127 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_2_zn 8.9fF
C128 comp_0_or3v0x2_0_zn comp_0_an3v0x2_1_a 4.1fF
C129 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_or2v0x3_0_zn 9.0fF
C130 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_2_zn 8.9fF
C131 totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_xor3v1x2_0_bn 2.6fF
C132 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_0_b 5.9fF
C133 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_an2v0x2_1_a 12.4fF
C134 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xor3v1x2_0_cn 18.8fF
C135 totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_0_mux_0_gnd 20.0fF
C136 totdiff3_0_mux_0_gnd comp_0_nr3v0x2_0_a 19.9fF
C137 totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_diff2_0_xor3v1x2_0_bn 2.4fF
C138 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xor3v1x2_0_cn 18.8fF
C139 totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_0_mux_0_gnd 9.1fF
C140 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_1_a 12.4fF
C141 totdiff3_0_mux_0_b2 totdiff3_0_mux_0_vdd 3.1fF
C142 totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_0_mux_0_mxn2v0x1_2_sn 9.2fF
C143 comp_0_an3v0x2_2_a comp_0_an3v0x2_0_zn 4.6fF
C144 comp_0_or3v0x2_1_zn totdiff3_0_mux_0_vdd 9.0fF
C145 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_in_b 4.3fF
C146 comp_0_an3v0x2_2_b totdiff3_0_mux_0_gnd 23.0fF
C147 comp_0_an3v0x2_2_w_n4_32# comp_0_an3v0x2_1_a 8.3fF
C148 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_bn 9.1fF
C149 totdiff3_0_mux_0_gnd comp_0_an3v0x2_3_zn 8.8fF
C150 comp_0_an3v0x2_2_a comp_0_iv1v0x4_2_a 2.2fF
C151 comp_0_an3v0x2_2_w_n4_32# comp_0_an3v0x2_2_z 21.1fF
C152 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_or2v0x3_0_zn 9.0fF
C153 comp_0_iv1v0x4_1_a totdiff3_0_mux_0_vdd 13.0fF
C154 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_diff2_2_xor2v2x2_0_bn 3.3fF
C155 totdiff3_1_diff2_0_an2v0x2_0_b totdiff3_0_mux_0_vdd 20.5fF
C156 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xor3v1x2_0_zn 11.9fF
C157 comp_0_or3v0x2_0_zn totdiff3_0_mux_0_gnd 10.9fF
C158 totdiff3_0_mux_0_a0 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 4.8fF
C159 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_a0 35.4fF
C160 totdiff3_1_mux_0_a2 totdiff3_0_mux_0_vdd 36.7fF
C161 comp_0_an3v0x2_2_a totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# 5.2fF
C162 totdiff3_1_mux_0_b1 totdiff3_1_diff2_1_xor2v2x2_0_bn 2.7fF
C163 totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_1_diff2_2_xor3v1x2_0_cn 2.3fF
C164 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xor2v2x2_0_an 27.4fF
C165 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_0_zn 10.8fF
C166 totdiff3_1_mux_0_s totdiff3_0_mux_0_gnd 8.3fF
C167 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_1_zn 8.9fF
C168 comp_0_an3v0x2_2_zn totdiff3_0_mux_0_vdd 4.9fF
C169 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_xor3v1x2_0_cn 18.8fF
C170 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_in_a 28.0fF
C171 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_s 36.4fF
C172 totdiff3_1_mux_0_b2 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 6.6fF
C173 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_1_a 20.0fF
C174 totdiff3_1_diff2_2_in_a totdiff3_0_mux_0_vdd 24.6fF
C175 totdiff3_1_diff2_1_an2v0x2_0_z totdiff3_0_mux_0_vdd 24.6fF
C176 comp_0_nd3v0x2_0_c totdiff3_0_mux_0_vdd 5.0fF
C177 totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 30.3fF
C178 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_s 7.9fF
C179 totdiff3_1_diff2_1_in_a totdiff3_1_diff2_1_an2v0x2_0_zn 2.2fF
C180 totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_diff2_1_xor2v2x2_0_an 3.3fF
C181 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_in_b 50.3fF
C182 totdiff3_0_mux_0_b2 totdiff3_0_mux_0_gnd 11.9fF
C183 totdiff3_1_mux_0_b0 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# 8.7fF
C184 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_1_a 20.0fF
C185 totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_mux_0_a1 4.1fF
C186 totdiff3_0_mux_0_gnd comp_0_or3v0x2_1_zn 10.9fF
C187 totdiff3_0_mux_0_gnd comp_0_iv1v0x4_1_a 8.9fF
C188 totdiff3_1_diff2_0_an2v0x2_0_b totdiff3_0_mux_0_gnd 7.3fF
C189 totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_xor3v1x2_0_zn 4.6fF
C190 comp_0_iv1v0x4_0_a totdiff3_0_mux_0_vdd 11.5fF
C191 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_a0 14.9fF
C192 totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_1_diff2_0_xor3v1x2_0_zn 4.5fF
C193 totdiff3_1_mux_0_b2 totdiff3_1_diff2_2_xor2v2x2_0_bn 2.7fF
C194 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_1_mux_0_b2 8.7fF
C195 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_1_mux_0_mxn2v0x1_2_zn 9.3fF
C196 totdiff3_1_mux_0_a2 totdiff3_0_mux_0_gnd 14.9fF
C197 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_xnr2v8x05_0_an 9.9fF
C198 totdiff3_0_mux_0_b0 totdiff3_0_diff2_0_xor2v2x2_0_an 3.9fF
C199 totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_1_diff2_0_xor3v1x2_0_cn 2.3fF
C200 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xor2v2x2_0_an 21.6fF
C201 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_diff2_0_xor3v1x2_0_cn 4.5fF
C202 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_vdd 59.4fF
C203 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_xor3v1x2_0_zn 18.9fF
C204 totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_xor3v1x2_0_zn 4.3fF
C205 totdiff3_1_diff2_2_an2v0x2_0_z totdiff3_0_mux_0_vdd 24.6fF
C206 comp_0_an3v0x2_2_zn totdiff3_0_mux_0_gnd 8.8fF
C207 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_mux_0_a2 4.1fF
C208 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_xnr2v8x05_0_zn 4.4fF
C209 totdiff3_0_diff2_2_an2v0x2_0_zn totdiff3_0_diff2_2_in_a 2.2fF
C210 totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_1_diff2_1_xor3v1x2_0_iz 2.4fF
C211 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_xnr2v8x05_0_zn 4.4fF
C212 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_1_mux_0_mxn2v0x1_0_zn 9.3fF
C213 totdiff3_0_mux_0_b2 totdiff3_0_diff2_2_xor2v2x2_0_bn 2.7fF
C214 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_1_mux_0_mxn2v0x1_2_zn 8.9fF
C215 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_vdd 18.9fF
C216 totdiff3_1_diff2_2_in_a totdiff3_0_mux_0_gnd 27.8fF
C217 totdiff3_1_diff2_1_an2v0x2_0_z totdiff3_0_mux_0_gnd 12.8fF
C218 comp_0_nd3v0x2_0_c totdiff3_0_mux_0_gnd 18.9fF
C219 totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_0_mux_0_vdd 17.7fF
C220 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_s 8.3fF
C221 totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_1_diff2_1_in_b 2.0fF
C222 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_in_b 60.8fF
C223 totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_0_mux_0_vdd 12.4fF
C224 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_xnr2v8x05_0_bn 14.4fF
C225 comp_0_an3v0x2_2_w_n4_32# comp_0_nr3v0x2_0_z 21.8fF
C226 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_1_zn 8.8fF
C227 totdiff3_1_diff2_1_in_c totdiff3_1_diff2_1_xnr2v8x05_0_zn 3.1fF
C228 comp_0_an3v0x2_2_w_n4_32# comp_0_nd3v0x2_0_a 6.2fF
C229 totdiff3_0_diff2_2_xnr2v8x05_0_an totdiff3_0_mux_0_vdd 9.9fF
C230 comp_0_iv1v0x4_0_a totdiff3_0_mux_0_gnd 11.2fF
C231 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_in_2c 33.2fF
C232 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xnr2v8x05_0_an 5.5fF
C233 totdiff3_1_mux_0_b0 totdiff3_0_mux_0_vdd 26.0fF
C234 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xor3v1x2_0_zn 18.9fF
C235 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xor3v1x2_0_zn 11.9fF
C236 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_xor3v1x2_0_cn 31.6fF
C237 totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_0_mux_0_vdd 12.7fF
C238 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_an2v0x2_0_z 12.8fF
C239 comp_0_an3v0x2_2_w_n4_32# comp_0_an3v0x2_0_z 9.5fF
C240 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_an2v0x2_1_z 17.9fF
C241 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xnr2v8x05_0_zn 15.0fF
C242 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xnr2v8x05_0_an 9.9fF
C243 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xnr2v8x05_0_zn 11.9fF
C244 comp_0_an3v0x2_2_a comp_0_an2v0x2_1_b 2.2fF
C245 totdiff3_0_mux_0_a0 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# 11.6fF
C246 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_gnd 11.9fF
C247 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_in_b 50.3fF
C248 totdiff3_0_diff2_2_an2v0x2_1_zn totdiff3_0_mux_0_vdd 8.8fF
C249 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_mxn2v0x1_2_zn 9.3fF
C250 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_xor2v2x2_0_bn 11.2fF
C251 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_0_mux_0_gnd 25.5fF
C252 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_xor3v1x2_0_cn 4.5fF
C253 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_an2v0x2_1_a 20.0fF
C254 totdiff3_1_diff2_2_in_c totdiff3_0_mux_0_vdd 40.7fF
C255 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xnr2v8x05_0_bn 6.7fF
C256 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_an2v0x2_1_z 17.9fF
C257 comp_0_an3v0x2_2_c totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# 6.3fF
C258 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_1_zn 8.9fF
C259 totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_1_diff2_0_xor3v1x2_0_bn 2.4fF
C260 totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_1_diff2_0_xor2v2x2_0_an 3.3fF
C261 totdiff3_1_diff2_2_in_c totdiff3_1_diff2_2_xnr2v8x05_0_zn 3.1fF
C262 totdiff3_1_diff2_2_in_b totdiff3_0_mux_0_vdd 50.3fF
C263 comp_0_an3v0x2_2_c comp_0_an3v0x2_0_b 2.7fF
C264 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xnr2v8x05_0_an 5.5fF
C265 totdiff3_0_mux_0_mxn2v0x1_0_sn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 9.2fF
C266 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_b1 6.6fF
C267 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_in_2c 17.8fF
C268 totdiff3_0_mux_0_b1 totdiff3_0_mux_0_a1 39.4fF
C269 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_or2v0x3_0_zn 12.7fF
C270 totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_diff2_1_xor2v2x2_0_bn 3.3fF
C271 comp_0_an3v0x2_2_c totdiff3_0_mux_0_vdd 25.3fF
C272 totdiff3_1_mux_0_b0 totdiff3_0_mux_0_gnd 10.9fF
C273 totdiff3_0_diff2_2_an2v0x2_2_z totdiff3_0_mux_0_vdd 2.4fF
C274 totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# 18.7fF
C275 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_zn 13.9fF
C276 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_cn 19.1fF
C277 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_1_mux_0_a1 13.4fF
C278 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_1_a 12.4fF
C279 totdiff3_0_mux_0_b1 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 10.2fF
C280 totdiff3_0_mux_0_b1 totdiff3_0_mux_0_vdd 13.1fF
C281 totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_0_mux_0_gnd 9.0fF
C282 totdiff3_1_diff2_2_an2v0x2_0_zn totdiff3_0_mux_0_vdd 8.8fF
C283 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_xor3v1x2_0_zn 18.9fF
C284 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_1_z 10.2fF
C285 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_an2v0x2_2_z 2.4fF
C286 totdiff3_0_mux_0_s totdiff3_0_mux_0_a2 4.5fF
C287 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xnr2v8x05_0_an 6.8fF
C288 totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_vdd 61.1fF
C289 totdiff3_1_diff2_1_an2v0x2_0_b totdiff3_0_mux_0_vdd 20.5fF
C290 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_1_mux_0_a0 11.6fF
C291 comp_0_iv1v0x4_2_a totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 5.0fF
C292 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_0_z 24.6fF
C293 comp_0_an2v0x2_0_b totdiff3_0_mux_0_vdd 49.9fF
C294 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xor3v1x2_0_cn 31.6fF
C295 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_in_b 60.8fF
C296 totdiff3_0_diff2_2_in_c totdiff3_0_mux_0_vdd 40.7fF
C297 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_1_zn 8.9fF
C298 comp_0_nd3v0x2_0_c comp_0_nr2v0x2_1_a 3.8fF
C299 comp_0_an3v0x2_2_w_n4_32# comp_0_nd3v0x2_0_z 5.2fF
C300 totdiff3_1_diff2_2_in_c totdiff3_0_mux_0_gnd 35.0fF
C301 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_an2v0x2_1_z 10.2fF
C302 totdiff3_1_mux_0_b1 totdiff3_1_diff2_1_xor2v2x2_0_an 3.9fF
C303 totdiff3_1_mux_0_b2 totdiff3_1_mux_0_mxn2v0x1_2_zn 2.7fF
C304 comp_0_an2v0x2_4_z totdiff3_0_mux_0_vdd 10.7fF
C305 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_in_b 60.5fF
C306 totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_xor3v1x2_0_zn 4.6fF
C307 totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_an2v0x2_1_a 2.0fF
C308 totdiff3_1_mux_0_b2 totdiff3_0_mux_0_vdd 3.1fF
C309 totdiff3_0_diff2_1_an2v0x2_2_zn totdiff3_0_mux_0_vdd 8.8fF
C310 comp_0_an3v0x2_1_a comp_0_an2v0x2_0_b 2.5fF
C311 comp_0_an3v0x2_2_c totdiff3_0_mux_0_gnd 36.3fF
C312 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_or2v0x3_0_zn 9.0fF
C313 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_a1 13.4fF
C314 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# comp_0_an3v0x2_0_b 5.0fF
C315 totdiff3_0_mux_0_b0 totdiff3_0_mux_0_b1 18.4fF
C316 totdiff3_0_diff2_2_an2v0x2_2_z totdiff3_0_mux_0_gnd 2.5fF
C317 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# 76.2fF
C318 totdiff3_0_mux_0_b1 totdiff3_0_mux_0_gnd 17.2fF
C319 totdiff3_1_diff2_2_an2v0x2_0_zn totdiff3_0_mux_0_gnd 8.9fF
C320 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_1_a 20.0fF
C321 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_vdd 59.4fF
C322 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_xor3v1x2_0_bn 15.4fF
C323 totdiff3_0_diff2_2_in_c totdiff3_0_diff2_2_xnr2v8x05_0_zn 3.1fF
C324 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_zn 13.9fF
C325 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_an2v0x2_2_z 2.5fF
C326 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_0_mux_0_a1 4.8fF
C327 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_a1 38.7fF
C328 comp_0_an3v0x2_0_b totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 2.3fF
C329 comp_0_an3v0x2_0_b totdiff3_0_mux_0_vdd 49.2fF
C330 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_an2v0x2_2_a 25.9fF
C331 totdiff3_1_diff2_1_an2v0x2_0_b totdiff3_0_mux_0_gnd 5.9fF
C332 totdiff3_1_mux_0_mxn2v0x1_1_zn totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 9.3fF
C333 comp_0_an2v0x2_0_b totdiff3_0_mux_0_gnd 32.8fF
C334 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_0_z 12.8fF
C335 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_cn 19.1fF
C336 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_in_b 50.3fF
C337 totdiff3_1_diff2_2_an2v0x2_1_z totdiff3_0_mux_0_vdd 17.9fF
C338 totdiff3_0_diff2_2_in_c totdiff3_0_mux_0_gnd 35.0fF
C339 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_an2v0x2_0_z 24.6fF
C340 totdiff3_1_diff2_2_xnr2v8x05_0_zn totdiff3_0_mux_0_vdd 4.4fF
C341 comp_0_an2v0x2_4_z totdiff3_0_mux_0_gnd 9.8fF
C342 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_an2v0x2_2_a 59.6fF
C343 totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_diff2_0_xor2v2x2_0_bn 3.3fF
C344 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_b2 11.9fF
C345 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_0_b 20.5fF
C346 totdiff3_1_diff2_1_in_c totdiff3_0_mux_0_vdd 39.6fF
C347 totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_0_mux_0_b2 8.7fF
C348 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_0_z 24.6fF
C349 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_2_zn 8.9fF
C350 comp_0_an3v0x2_1_a totdiff3_0_mux_0_vdd 72.4fF
C351 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_1_mux_0_a1 4.8fF
C352 comp_0_an3v0x2_2_z totdiff3_0_mux_0_vdd 3.3fF
C353 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_xnr2v8x05_0_bn 14.4fF
C354 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_xnr2v8x05_0_zn 4.4fF
C355 totdiff3_0_mux_0_mxn2v0x1_0_zn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 8.9fF
C356 comp_0_an3v0x2_2_a comp_0_or3v0x2_0_zn 3.3fF
C357 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xor3v1x2_0_bn 9.1fF
C358 comp_0_iv1v0x4_1_a totdiff3_1_mux_0_a0 2.3fF
C359 totdiff3_1_diff2_0_an2v0x2_0_zn totdiff3_0_mux_0_vdd 8.8fF
C360 totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_1_diff2_1_xor3v1x2_0_cn 2.3fF
C361 totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_vdd 59.6fF
C362 totdiff3_0_diff2_0_an2v0x2_0_b totdiff3_0_mux_0_vdd 20.5fF
C363 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# comp_0_iv1v0x4_2_a 2.3fF
C364 comp_0_an3v0x2_0_b totdiff3_0_mux_0_gnd 34.1fF
C365 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_an2v0x2_1_z 17.9fF
C366 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_a1 15.3fF
C367 totdiff3_0_mux_0_b0 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 8.7fF
C368 totdiff3_0_mux_0_b0 totdiff3_0_mux_0_vdd 26.0fF
C369 totdiff3_0_mux_0_mxn2v0x1_0_sn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# 9.3fF
C370 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_in_b 60.5fF
C371 totdiff3_1_diff2_2_an2v0x2_1_z totdiff3_0_mux_0_gnd 10.2fF
C372 totdiff3_1_mux_0_b0 totdiff3_1_mux_0_mxn2v0x1_0_zn 2.7fF
C373 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_vdd 92.6fF
C374 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 76.0fF
C375 comp_0_an3v0x2_2_a comp_0_an3v0x2_2_w_n4_32# 8.7fF
C376 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_in_a 24.6fF
C377 totdiff3_0_diff2_1_an2v0x2_1_a totdiff3_0_diff2_1_in_b 2.0fF
C378 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_0_z 12.8fF
C379 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_xnr2v8x05_0_zn 11.9fF
C380 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_2_a 59.6fF
C381 comp_0_an2v0x2_3_z totdiff3_0_mux_0_vdd 9.1fF
C382 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_an2v0x2_2_a 25.9fF
C383 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xnr2v8x05_0_bn 14.4fF
C384 comp_0_an3v0x2_2_w_n4_32# comp_0_an3v0x2_1_zn 5.8fF
C385 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_0_b 5.9fF
C386 totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_0_mux_0_s 15.2fF
C387 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_an2v0x2_1_a 12.4fF
C388 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_in_c 34.1fF
C389 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_0_z 12.8fF
C390 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_1_mux_0_s 18.7fF
C391 totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_an2v0x2_1_a 2.0fF
C392 totdiff3_1_diff2_2_an2v0x2_2_zn totdiff3_0_mux_0_vdd 8.8fF
C393 totdiff3_0_mux_0_mxn2v0x1_0_zn totdiff3_0_mux_0_b0 2.7fF
C394 comp_0_an3v0x2_1_a totdiff3_0_mux_0_gnd 57.3fF
C395 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xnr2v8x05_0_bn 6.7fF
C396 comp_0_an3v0x2_2_z totdiff3_0_mux_0_gnd 10.7fF
C397 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xnr2v8x05_0_zn 11.9fF
C398 totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_diff2_0_in_b 2.6fF
C399 comp_0_an2v0x2_2_z totdiff3_0_mux_0_vdd 9.4fF
C400 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_xor2v2x2_0_bn 17.7fF
C401 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_an2v0x2_0_zn 10.8fF
C402 totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_gnd 25.9fF
C403 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_0_b 7.3fF
C404 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_an2v0x2_1_z 10.2fF
C405 comp_0_an3v0x2_2_a totdiff3_0_mux_0_a0 2.3fF
C406 totdiff3_1_diff2_2_xnr2v8x05_0_bn totdiff3_0_mux_0_vdd 14.4fF
C407 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_an2v0x2_0_zn 8.8fF
C408 totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_diff2_1_xor3v1x2_0_zn 4.5fF
C409 totdiff3_1_mux_0_mxn2v0x1_1_zn totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# 8.9fF
C410 totdiff3_0_mux_0_b0 totdiff3_0_mux_0_gnd 10.9fF
C411 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_xor3v1x2_0_bn 15.4fF
C412 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_1_mux_0_mxn2v0x1_0_zn 8.9fF
C413 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_a1 38.7fF
C414 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_in_a 27.8fF
C415 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# comp_0_iv1v0x4_1_a 5.2fF
C416 comp_0_an3v0x2_2_w_n4_32# comp_0_nr3v0x2_0_a 15.0fF
C417 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_2_a 25.9fF
C418 totdiff3_0_mux_0_b2 totdiff3_0_diff2_2_xor2v2x2_0_an 3.9fF
C419 comp_0_an3v0x2_0_zn totdiff3_0_mux_0_vdd 10.7fF
C420 totdiff3_0_diff2_1_xor3v1x2_0_bn totdiff3_0_diff2_1_in_b 2.6fF
C421 comp_0_an2v0x2_3_z totdiff3_0_mux_0_gnd 20.8fF
C422 comp_0_an2v0x2_0_zn totdiff3_0_mux_0_vdd 8.8fF
C423 comp_0_an3v0x2_2_w_n4_32# comp_0_an3v0x2_2_b 21.4fF
C424 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_xnr2v8x05_0_bn 14.4fF
C425 comp_0_iv1v0x4_2_a totdiff3_0_mux_0_vdd 13.7fF
C426 totdiff3_1_mux_0_mxn2v0x1_2_sn totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 9.3fF
C427 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xnr2v8x05_0_bn 7.5fF
C428 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_xor3v1x2_0_iz 15.8fF
C429 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_in_b 50.3fF
C430 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_an2v0x2_1_a 20.0fF
C431 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_a2 11.6fF
C432 totdiff3_1_diff2_1_an2v0x2_2_zn totdiff3_0_mux_0_vdd 8.8fF
C433 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_xnr2v8x05_0_an 9.9fF
C434 totdiff3_1_diff2_2_an2v0x2_2_zn totdiff3_0_mux_0_gnd 8.9fF
C435 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# 21.1fF
C436 totdiff3_1_diff2_2_in_2c totdiff3_0_mux_0_vdd 33.2fF
C437 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_diff2_2_xor2v2x2_0_bn 3.3fF
C438 comp_0_nr3v0x2_0_z totdiff3_0_mux_0_vdd 8.7fF
C439 totdiff3_1_mux_0_b1 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 6.6fF
C440 comp_0_nd3v0x2_0_a totdiff3_0_mux_0_vdd 9.6fF
C441 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_an2v0x2_0_b 20.5fF
C442 totdiff3_0_mux_0_vdd totdiff3_0_mux_0_a2 36.7fF
C443 totdiff3_1_mux_0_b0 totdiff3_1_diff2_0_xor2v2x2_0_bn 2.7fF
C444 totdiff3_0_mux_0_gnd comp_0_an2v0x2_2_z 11.1fF
C445 comp_0_an3v0x2_1_a comp_0_an3v0x2_0_zn 2.5fF
C446 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xor2v2x2_0_bn 11.2fF
C447 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_xor3v1x2_0_iz 15.8fF
C448 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_1_mux_0_mxn2v0x1_2_sn 9.2fF
C449 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_mxn2v0x1_1_sn 9.3fF
C450 totdiff3_0_diff2_0_an2v0x2_0_zn totdiff3_0_diff2_0_in_a 2.2fF
C451 totdiff3_1_diff2_2_xnr2v8x05_0_bn totdiff3_0_mux_0_gnd 6.7fF
C452 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_xnr2v8x05_0_zn 4.4fF
C453 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_an2v0x2_0_zn 8.9fF
C454 totdiff3_0_diff2_1_an2v0x2_0_zn totdiff3_0_diff2_1_in_a 2.2fF
C455 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xor3v1x2_0_iz 15.8fF
C456 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xor3v1x2_0_bn 9.1fF
C457 totdiff3_0_mux_0_vdd totdiff3_1_diff2_1_xor2v2x2_0_bn 17.7fF
C458 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_mxn2v0x1_2_sn 9.3fF
C459 totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_diff2_1_xor3v1x2_0_bn 2.4fF
C460 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_1_mux_0_mxn2v0x1_0_sn 9.3fF
C461 totdiff3_0_mux_0_gnd totdiff3_1_mux_0_a1 15.3fF
C462 comp_0_nr2v0x2_1_a totdiff3_0_mux_0_vdd 7.1fF
C463 totdiff3_0_mux_0_mxn2v0x1_1_sn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 9.2fF
C464 totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_xor3v1x2_0_bn 2.6fF
C465 totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_1_mux_0_a0 4.1fF
C466 totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_xor3v1x2_0_zn 4.3fF
C467 totdiff3_0_mux_0_gnd comp_0_an3v0x2_0_zn 8.8fF
C468 comp_0_an3v0x2_0_z totdiff3_0_mux_0_vdd 2.3fF
C469 totdiff3_0_mux_0_mxn2v0x1_0_zn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# 9.3fF
C470 totdiff3_0_mux_0_gnd comp_0_an2v0x2_0_zn 8.9fF
C471 comp_0_an3v0x2_2_zn comp_0_nr3v0x2_0_a 2.1fF
C472 totdiff3_0_mux_0_gnd comp_0_iv1v0x4_2_a 9.0fF
C473 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_in_a 24.6fF
C474 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xnr2v8x05_0_bn 6.7fF
C475 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_xor3v1x2_0_iz 15.8fF
C476 totdiff3_0_mux_0_gnd totdiff3_0_diff2_2_xor3v1x2_0_iz 24.9fF
C477 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_in_b 60.5fF
C478 totdiff3_0_mux_0_b0 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# 6.6fF
C479 totdiff3_1_mux_0_mxn2v0x1_1_sn totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 9.3fF
C480 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_xnr2v8x05_0_bn 14.4fF
C481 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xnr2v8x05_0_an 5.5fF
C482 totdiff3_1_diff2_1_an2v0x2_2_zn totdiff3_0_mux_0_gnd 8.9fF
C483 totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_0_mux_0_vdd 15.8fF
C484 totdiff3_1_mux_0_s totdiff3_1_mux_0_a2 4.5fF
C485 totdiff3_1_diff2_2_in_2c totdiff3_0_mux_0_gnd 17.8fF
C486 totdiff3_1_mux_0_b0 totdiff3_1_mux_0_b1 18.4fF
C487 comp_0_nr3v0x2_0_z totdiff3_0_mux_0_gnd 21.2fF
C488 totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_xor3v1x2_0_cn 4.1fF
C489 comp_0_nd3v0x2_0_a totdiff3_0_mux_0_gnd 21.1fF
C490 totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_0_mux_0_mxn2v0x1_2_zn 8.9fF
C491 totdiff3_0_mux_0_gnd totdiff3_1_diff2_2_an2v0x2_0_b 5.9fF
C492 comp_0_an2v0x2_4_zn totdiff3_0_mux_0_vdd 8.8fF
C493 totdiff3_0_mux_0_gnd totdiff3_0_mux_0_a2 14.9fF
C494 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xor3v1x2_0_iz 24.9fF
C495 totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# comp_0_an3v0x2_2_c 2.3fF
C496 totdiff3_0_mux_0_vdd comp_0_an2v0x2_2_zn 8.8fF
C497 comp_0_an3v0x2_2_w_n4_32# comp_0_an3v0x2_2_zn 5.8fF
C498 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xnr2v8x05_0_zn 11.9fF
C499 totdiff3_0_mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_iz 25.5fF
C500 totdiff3_0_mux_0_gnd totdiff3_1_diff2_1_xor2v2x2_0_bn 11.2fF
C501 totdiff3_1_diff2_1_in_a totdiff3_0_mux_0_vdd 24.6fF
C502 totdiff3_0_mux_0_b1 totdiff3_0_diff2_1_xor2v2x2_0_an 3.9fF
C503 totdiff3_1_diff2_0_an2v0x2_0_zn totdiff3_1_diff2_0_in_a 2.2fF
C504 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_xor3v1x2_0_iz 15.8fF
C505 totdiff3_1_mux_0_b0 totdiff3_1_diff2_0_xor2v2x2_0_an 3.9fF
C506 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_1_mux_0_a0 4.8fF
C507 comp_0_nr2v0x2_1_a totdiff3_0_mux_0_gnd 22.9fF
C508 comp_0_nd3v0x2_0_c comp_0_an3v0x2_2_w_n4_32# 5.7fF
C509 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_xor3v1x2_0_zn 4.5fF
C510 comp_0_an3v0x2_0_z totdiff3_0_mux_0_gnd 36.9fF
C511 totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_xor3v1x2_0_zn 4.6fF
C512 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_in_a 28.0fF
C513 totdiff3_0_mux_0_gnd totdiff3_0_diff2_1_xor3v1x2_0_iz 24.9fF
C514 totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_diff2_2_xor3v1x2_0_bn 2.4fF
C515 comp_0_an2v0x2_3_b totdiff3_0_mux_0_vdd 13.7fF
C516 totdiff3_1_mux_0_b0 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# 6.6fF
C517 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xnr2v8x05_0_bn 7.5fF
C518 totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_0_mux_0_gnd 24.9fF
C519 comp_0_nd3v0x2_0_z totdiff3_0_mux_0_vdd 6.1fF
C520 comp_0_an3v0x2_2_a totdiff3_1_diff2_2_in_c 9.3fF
C521 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_in_c 39.6fF
C522 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_1_mux_0_b1 10.2fF
C523 totdiff3_0_mux_0_vdd totdiff3_0_diff2_0_xor2v2x2_0_bn 18.7fF
C524 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_an2v0x2_1_zn 8.8fF
C525 totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 36.4fF
C526 totdiff3_0_mux_0_gnd comp_0_an2v0x2_4_zn 8.9fF
C527 totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_diff2_0_in_b 2.0fF
C528 totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_diff2_0_xor3v1x2_0_cn 2.3fF
C529 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_an2v0x2_0_zn 8.8fF
C530 totdiff3_0_mux_0_gnd comp_0_an2v0x2_2_zn 8.9fF
C531 comp_0_an3v0x2_2_a totdiff3_0_mux_0_mxn2v0x1_0_sn 4.3fF
C532 totdiff3_0_mux_0_vdd totdiff3_1_diff2_2_xor3v1x2_0_bn 15.4fF
C533 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_mux_0_b2 3.9fF
C534 comp_0_an2v0x2_1_b totdiff3_0_mux_0_vdd 14.2fF
C535 totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_xor3v1x2_0_zn 4.6fF
C536 totdiff3_1_mux_0_mxn2v0x1_0_sn comp_0_iv1v0x4_1_a 4.3fF
C537 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_or2v0x3_0_zn 12.7fF
C538 totdiff3_1_diff2_1_in_a totdiff3_0_mux_0_gnd 27.8fF
C539 totdiff3_0_mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_iz 25.5fF
C540 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_1_mux_0_s 15.2fF
C541 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_xor3v1x2_0_zn 18.9fF
C542 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_xor3v1x2_0_cn 4.5fF
C543 totdiff3_0_mux_0_vdd totdiff3_1_diff2_0_xor2v2x2_0_bn 18.7fF
C544 comp_0_an2v0x2_3_b totdiff3_0_mux_0_gnd 15.0fF
C545 totdiff3_0_mux_0_b1 totdiff3_0_diff2_1_xor2v2x2_0_bn 2.7fF
C546 comp_0_an3v0x2_2_a comp_0_an2v0x2_0_b 4.9fF
C547 totdiff3_0_mux_0_vdd totdiff3_0_diff2_1_xor2v2x2_0_an 25.5fF
C548 totdiff3_1_mux_0_mxn2v0x1_1_sn totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# 9.2fF
C549 totdiff3_0_mux_0_vdd totdiff3_1_mux_0_a0 35.4fF
C550 totdiff3_1_mux_0_a2 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 11.6fF
C551 totdiff3_1_diff2_0_an2v0x2_2_zn totdiff3_0_mux_0_vdd 10.3fF
C552 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_vdd 25.5fF
C553 comp_0_nd3v0x2_0_z totdiff3_0_mux_0_gnd 5.3fF
C554 totdiff3_0_mux_0_vdd totdiff3_0_diff2_2_in_a 24.6fF
C555 totdiff3_0_mux_0_b0 totdiff3_0_diff2_0_xor2v2x2_0_bn 2.7fF
C556 totdiff3_1_diff2_1_an2v0x2_0_zn totdiff3_0_mux_0_vdd 8.8fF
C557 totdiff3_0_diff2_0_in_a 0 4.4fF
C558 totdiff3_0_diff2_0_an2v0x2_0_b 0 2.9fF
C559 totdiff3_0_diff2_1_in_c 0 37.1fF
C560 totdiff3_0_diff2_0_an2v0x2_0_z 0 5.0fF
C561 totdiff3_0_diff2_1_in_a 0 4.4fF
C562 totdiff3_0_mux_0_a1 0 28.9fF
C563 totdiff3_0_diff2_1_an2v0x2_0_b 0 2.9fF
C564 totdiff3_0_diff2_2_in_c 0 36.8fF
C565 totdiff3_0_diff2_1_an2v0x2_0_z 0 5.0fF
C566 totdiff3_0_diff2_1_in_2c 0 29.6fF
C567 totdiff3_0_diff2_2_in_a 0 4.4fF
C568 totdiff3_0_mux_0_a2 0 38.7fF
C569 totdiff3_0_diff2_2_an2v0x2_0_b 0 2.9fF
C570 totdiff3_0_diff2_2_an2v0x2_0_z 0 5.0fF
C571 totdiff3_0_diff2_2_in_2c 0 34.8fF
C572 comp_0_an3v0x2_2_a 0 184.1fF
C573 totdiff3_0_mux_0_b0 0 47.5fF
C574 totdiff3_0_mux_0_s 0 16.3fF
C575 totdiff3_0_mux_0_a0 0 99.1fF
C576 totdiff3_0_mux_0_b1 0 87.1fF
C577 totdiff3_0_mux_0_b2 0 24.6fF
C578 totdiff3_1_diff2_0_in_a 0 4.4fF
C579 totdiff3_1_diff2_0_an2v0x2_0_b 0 2.9fF
C580 totdiff3_1_diff2_1_in_c 0 37.1fF
C581 totdiff3_1_diff2_0_an2v0x2_0_z 0 5.0fF
C582 totdiff3_1_diff2_1_in_a 0 4.4fF
C583 totdiff3_1_mux_0_a1 0 28.9fF
C584 totdiff3_1_diff2_1_an2v0x2_0_b 0 2.9fF
C585 totdiff3_1_diff2_2_in_c 0 36.8fF
C586 totdiff3_1_diff2_1_an2v0x2_0_z 0 5.0fF
C587 totdiff3_1_diff2_1_in_2c 0 29.6fF
C588 totdiff3_1_diff2_2_in_a 0 4.4fF
C589 totdiff3_1_mux_0_a2 0 38.7fF
C590 totdiff3_1_diff2_2_an2v0x2_0_b 0 2.9fF
C591 totdiff3_1_diff2_2_an2v0x2_0_z 0 5.0fF
C592 totdiff3_1_diff2_2_in_2c 0 34.8fF
C593 totdiff3_1_mux_0_b0 0 47.5fF
C594 totdiff3_1_mux_0_s 0 16.3fF
C595 totdiff3_1_mux_0_a0 0 99.1fF
C596 totdiff3_1_mux_0_b1 0 87.1fF
C597 totdiff3_1_mux_0_b2 0 24.6fF
C598 comp_0_iv1v0x4_0_a 0 24.2fF
C599 comp_0_iv1v0x4_1_a 0 15.1fF
C600 comp_0_an3v0x2_0_b 0 78.6fF
C601 comp_0_an3v0x2_2_c 0 98.7fF
C602 totdiff3_0_mux_0_vdd 0 663.6fF
C603 comp_0_iv1v0x4_2_a 0 19.0fF
C604 totdiff3_0_mux_0_gnd 0 794.7fF
C605 comp_0_nr3v0x2_0_a 0 8.6fF

v_dd totdiff3_0_mux_0_vdd 0 5
v_ss totdiff3_0_mux_0_gnd 0 0

v_a11 totdiff3_0_diff2_0_in_a 0 DC 1 PULSE(0 5 0 0 0 20ns 40ns )
v_a12 totdiff3_0_diff2_1_in_a 0 DC 1 PULSE(0 5 0 0 0 20ns 40ns )
v_a13 totdiff3_0_diff2_2_in_a 0 DC 1 PULSE(0 5 0 0 0 20ns 40ns )
v_b11 totdiff3_0_diff2_0_in_b 0 DC 1 PULSE(0 5 0 0 0 40ns 80ns )
v_b12 totdiff3_0_diff2_1_in_b 0 DC 1 PULSE(0 5 0 0 0 40ns 80ns )
v_b13 totdiff3_0_diff2_2_in_b 0 DC 1 PULSE(0 5 0 0 0 40ns 80ns )


v_a21 totdiff3_1_diff2_0_in_a 0 DC 1 PULSE(0 5 0 0 0 20ns 40ns )
v_a22 totdiff3_1_diff2_1_in_a 0 DC 1 PULSE(0 5 0 0 0 20ns 40ns )
v_a23 totdiff3_1_diff2_2_in_a 0 DC 1 PULSE(0 5 0 0 0 20ns 40ns )
v_b21 totdiff3_1_diff2_0_in_b 0 DC 1 PULSE(0 5 0 0 0 40ns 80ns )
v_b22 totdiff3_1_diff2_1_in_b 0 DC 1 PULSE(0 5 0 0 0 40ns 80ns )
v_b23 totdiff3_1_diff2_2_in_b 0 DC 1 PULSE(0 5 0 0 0 40ns 80ns )

.tran 0.1ns 200ns 
comp_0_iv1v0x4_0_a
.control
run 
setplot tran1
plot comp_0_nd3v0x2_0_z
.endc 

.end