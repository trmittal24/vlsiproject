* Mon Aug 16 14:22:56 CEST 2004
.subckt inv_x4 i nq vdd vss 
*SPICE circuit <inv_x4> from XCircuit v3.10

m1 nq i vss vss n w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m2 nq i vdd vdd p w=68u l=2u ad='68u*5u+12p' as='68u*5u+12p' pd='68u*2+14u' ps='68u*2+14u'
.ends
