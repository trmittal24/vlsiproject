* Spice description of oai21_x05
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:10
*
.subckt oai21_x05 a1 a2 b vdd vss z 
M3  vdd   b     z     vdd p  L=0.13U  W=0.605U AS=0.160325P AD=0.160325P PS=1.74U   PD=1.74U  
M2  z     a2    n1    vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M1  n1    a1    vdd   vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M6  n2    b     z     vss n  L=0.13U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U  
M5  vss   a2    n2    vss n  L=0.13U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U  
M4  n2    a1    vss   vss n  L=0.13U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U  
C8  a1    vss   1.067f
C7  b     vss   1.410f
C6  a2    vss   1.056f
C4  vdd   vss   1.114f
C3  z     vss   2.163f
C2  n2    vss   0.529f
.ends
