* Sat Aug 27 19:34:25 CEST 2005
.subckt nd2v4x1 a b vdd vss z 
*SPICE circuit <nd2v4x1> from XCircuit v3.20

m1 n1 a vss vss n w=8u l=2.3636u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
m2 z a vdd vdd p w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m3 z b n1 vss n w=8u l=2.3636u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
m4 z b vdd vdd p w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
.ends
