* Sat Mar 31 18:39:50 CEST 2007
.subckt nd2v6x3 a b vdd vss z
*SPICE circuit <nd2v6x3> from XCircuit v3.4 rev 26

m1 n1 a vss vss n w=30u l=2.3636u ad='30u*5u+12p' as='30u*5u+12p' pd='30u*2+14u' ps='30u*2+14u'
m2 z a vdd vdd p w=36u l=2.3636u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
m3 z b n1 vss n w=30u l=2.3636u ad='30u*5u+12p' as='30u*5u+12p' pd='30u*2+14u' ps='30u*2+14u'
m4 z b vdd vdd p w=36u l=2.3636u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
.ends
