* Mon Aug 16 14:22:57 CEST 2004
.subckt o3_x2 i0 i1 i2 q vdd vss 
*SPICE circuit <o3_x2> from XCircuit v3.10

m1 nq i2 n2 vdd p w=30u l=2.3636u ad='30u*5u+12p' as='30u*5u+12p' pd='30u*2+14u' ps='30u*2+14u'
m2 n2 i1 n1 vdd p w=30u l=2.3636u ad='30u*5u+12p' as='30u*5u+12p' pd='30u*2+14u' ps='30u*2+14u'
m3 q nq vdd vdd p w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m4 q nq vss vss n w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m5 nq i0 vss vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m6 nq i1 vss vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m7 nq i2 vss vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m8 n1 i0 vdd vdd p w=30u l=2.3636u ad='30u*5u+12p' as='30u*5u+12p' pd='30u*2+14u' ps='30u*2+14u'
.ends
