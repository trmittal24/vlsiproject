* Spice description of nd3_x2
* Spice driver version 134999461
* Date 31/05/2007 at 21:34:33
* vxlib 0.13um values
.subckt nd3_x2 a b c vdd vss z
M1a z     a     vdd   vdd p  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M1b vdd   b     z     vdd p  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M1z z     c     vdd   vdd p  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M2a vss   a     sig1  vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M2b sig1  b     n2    vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M2c n2    c     z     vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
C7  a     vss   0.749f
C6  b     vss   0.655f
C8  c     vss   0.533f
C4  z     vss   1.287f
.ends
