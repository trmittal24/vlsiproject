* Spice description of nd2av0x05
* Spice driver version 134999461
* Date 17/05/2007 at  9:16:58
* vsclib 0.13um values
.subckt nd2av0x05 a b vdd vss z
M01 06    a     vdd   vdd p  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
M02 06    a     vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M03 z     b     vdd   vdd p  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M04 sig3  b     z     vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M05 vdd   06    z     vdd p  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M06 vss   06    sig3  vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
C5  06    vss   0.559f
C6  a     vss   0.476f
C4  b     vss   0.506f
C2  z     vss   0.513f
.ends
