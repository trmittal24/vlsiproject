* Sat Apr  9 11:25:46 CEST 2005
.subckt nr2v0x8 a b vdd vss z 
*SPICE circuit <nr2v0x8> from XCircuit v3.20

m1 z a vss vss n w=58u l=2u ad='58u*5u+12p' as='58u*5u+12p' pd='58u*2+14u' ps='58u*2+14u'
m2 n1 a vdd vdd p w=216u l=2u ad='216u*5u+12p' as='216u*5u+12p' pd='216u*2+14u' ps='216u*2+14u'
m3 z b vss vss n w=58u l=2u ad='58u*5u+12p' as='58u*5u+12p' pd='58u*2+14u' ps='58u*2+14u'
m4 z b n1 vdd p w=216u l=2u ad='216u*5u+12p' as='216u*5u+12p' pd='216u*2+14u' ps='216u*2+14u'
.ends
