* Spice description of nd4_x05
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:10
*
.subckt nd4_x05 a b c d vdd vss z 
M4  vdd   a     z     vdd p  L=0.13U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U  
M3  z     b     vdd   vdd p  L=0.13U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U  
M2  vdd   c     z     vdd p  L=0.13U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U  
M1  z     d     vdd   vdd p  L=0.13U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U  
M8  sig2  a     vss   vss n  L=0.13U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U  
M7  sig1  b     sig2  vss n  L=0.13U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U  
M5  z     d     n3    vss n  L=0.13U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U  
M6  n3    c     sig1  vss n  L=0.13U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U  
C10 vdd   vss   1.860f
C9  b     vss   1.002f
C8  d     vss   1.035f
C7  c     vss   0.767f
C6  a     vss   0.989f
C4  z     vss   2.574f
.ends
