* Fri May  4 21:00:20 CEST 2007
.subckt xnai21v0x05 a1 a2 b vdd vss z
*SPICE circuit <xnai21v0x05> from XCircuit v3.4 rev 26

m1 z b vdd vdd p w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m2 n2 b vss vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m3 z a2n a1n vdd p w=21u l=2.3636u ad='21u*5u+12p' as='21u*5u+12p' pd='21u*2+14u' ps='21u*2+14u'
m4 a2n a2 vss vss n w=11u l=2.3636u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m5 a1n a1 n2 vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m6 z a1n n1 vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m7 n1 a2n n2 vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m8 a1n a1 vdd vdd p w=21u l=2.3636u ad='21u*5u+12p' as='21u*5u+12p' pd='21u*2+14u' ps='21u*2+14u'
m9 a2n a2 vdd vdd p w=21u l=2.3636u ad='21u*5u+12p' as='21u*5u+12p' pd='21u*2+14u' ps='21u*2+14u'
m10 z a2 a1n vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m11 z a1n a2n vdd p w=21u l=2.3636u ad='21u*5u+12p' as='21u*5u+12p' pd='21u*2+14u' ps='21u*2+14u'
.ends
