* Spice description of nd2v0x2
* Spice driver version 134894944
* Date  4/10/2005 at 10:05:30
*
.subckt nd2v0x2 a b vdd vss z 
M1b z     b     vdd   vdd p  L=0.12U  W=1.32U  AS=0.363P    AD=0.363P    PS=3.19U   PD=3.19U  
M1a vdd   a     z     vdd p  L=0.12U  W=1.32U  AS=0.363P    AD=0.363P    PS=3.19U   PD=3.19U  
M2b n1    b     z     vss n  L=0.12U  W=1.1U   AS=0.3025P   AD=0.3025P   PS=2.75U   PD=2.75U  
M2a vss   a     n1    vss n  L=0.12U  W=1.1U   AS=0.3025P   AD=0.3025P   PS=2.75U   PD=2.75U  
C6  vdd   vss   0.808f
C5  b     vss   0.468f
C4  a     vss   0.600f
C3  z     vss   0.499f
.ends
