* Spice description of nd2v5x1
* Spice driver version 134999461
* Date 17/05/2007 at  9:20:52
* wsclib 0.13um values
.subckt nd2v5x1 a b vdd vss z
M01 vdd   a     z     vdd p  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
M02 vss   a     n1    vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M03 z     b     vdd   vdd p  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
M04 n1    b     z     vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
C4  a     vss   0.409f
C5  b     vss   0.353f
C1  z     vss   0.674f
.ends
