* Tue Aug 10 11:21:07 CEST 2004
.subckt nd4_x2 a b c d vdd vss z 
*SPICE circuit <nd4_x2> from XCircuit v3.10

m1 n1 a vss vss n w=46u l=2u ad='46u*5u+12p' as='46u*5u+12p' pd='46u*2+14u' ps='46u*2+14u'
m2 n2 b n1 vss n w=46u l=2u ad='46u*5u+12p' as='46u*5u+12p' pd='46u*2+14u' ps='46u*2+14u'
m3 n3 c n2 vss n w=46u l=2u ad='46u*5u+12p' as='46u*5u+12p' pd='46u*2+14u' ps='46u*2+14u'
m4 z d n3 vss n w=46u l=2u ad='46u*5u+12p' as='46u*5u+12p' pd='46u*2+14u' ps='46u*2+14u'
m5 z a vdd vdd p w=39u l=2u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m6 z b vdd vdd p w=39u l=2u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m7 z c vdd vdd p w=39u l=2u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m8 z d vdd vdd p w=39u l=2u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
.ends
