* Spice description of nd3_x05
* Spice driver version 134999461
* Date 31/05/2007 at 21:34:29
* vxlib 0.13um values
.subckt nd3_x05 a b c vdd vss z
M1  z     c     vdd   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M2  vdd   b     z     vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M3  z     a     vdd   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M4  sig4  c     z     vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M5  n1    b     sig4  vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M6  vss   a     n1    vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
C5  a     vss   0.610f
C7  b     vss   0.594f
C6  c     vss   0.604f
C3  z     vss   1.040f
.ends
