* Fri Apr  8 11:37:18 CEST 2005
.subckt aoi31v0x3 a1 a2 a3 b vdd vss z 
*SPICE circuit <aoi31v0x3> from XCircuit v3.20

m1 n1 a1 vss vss n w=54u l=2u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m2 n3 a1 vdd vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m3 n3 a3 vdd vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m4 n3 a2 vdd vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m5 n2 a2 n1 vss n w=54u l=2u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m6 z b vss vss n w=22u l=2u ad='22u*5u+12p' as='22u*5u+12p' pd='22u*2+14u' ps='22u*2+14u'
m7 z a3 n2 vss n w=54u l=2u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m8 z b n3 vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
.ends
