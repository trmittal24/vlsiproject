* Sat Apr  9 10:46:05 CEST 2005
.subckt nd2av0x6 a b vdd vss z 
*SPICE circuit <nd2av0x6> from XCircuit v3.20

m1 an a vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m2 n1 b vss vss n w=60u l=2u ad='60u*5u+12p' as='60u*5u+12p' pd='60u*2+14u' ps='60u*2+14u'
m3 an a vdd vdd p w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m4 z b vdd vdd p w=72u l=2u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
m5 z an n1 vss n w=60u l=2u ad='60u*5u+12p' as='60u*5u+12p' pd='60u*2+14u' ps='60u*2+14u'
m6 z an vdd vdd p w=72u l=2u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
.ends
