* Tue Feb 20 08:57:11 CET 2007
.subckt nr2av0x1 a b vdd vss z
*SPICE circuit <nr2av0x1> from XCircuit v3.4 rev 26

m1 an a vss vss n w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m2 an a vdd vdd p w=26u l=2.3636u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m3 z an vss vss n w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m4 n1 an vdd vdd p w=26u l=2.3636u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m5 z b vss vss n w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m6 z b n1 vdd p w=26u l=2.3636u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
.ends
