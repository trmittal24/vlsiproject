* Sun Apr  2 21:56:05 CEST 2006
.subckt nd2v3x4 a b vdd vss z 
*SPICE circuit <nd2v3x4> from XCircuit v3.20

m1 n1 a vss vss n w=80u l=2.3636u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m2 z a vdd vdd p w=48u l=2.3636u ad='48u*5u+12p' as='48u*5u+12p' pd='48u*2+14u' ps='48u*2+14u'
m3 z b n1 vss n w=80u l=2.3636u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m4 z b vdd vdd p w=48u l=2.3636u ad='48u*5u+12p' as='48u*5u+12p' pd='48u*2+14u' ps='48u*2+14u'
.ends
