* Wed May  2 18:42:06 CEST 2007
.subckt mxi2v2x3 a0 a1 s vdd vss z
*SPICE circuit <mxi2v2x3> from XCircuit v3.4 rev 26

m1 a0n a0 vdd vdd p w=66u l=2.3636u ad='66u*5u+12p' as='66u*5u+12p' pd='66u*2+14u' ps='66u*2+14u'
m2 a1n a1 vdd vdd p w=66u l=2.3636u ad='66u*5u+12p' as='66u*5u+12p' pd='66u*2+14u' ps='66u*2+14u'
m3 z sn a1n vdd p w=66u l=2.3636u ad='66u*5u+12p' as='66u*5u+12p' pd='66u*2+14u' ps='66u*2+14u'
m4 a0n s z vdd p w=66u l=2.3636u ad='66u*5u+12p' as='66u*5u+12p' pd='66u*2+14u' ps='66u*2+14u'
m5 sn s vdd vdd p w=24u l=2.3636u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m6 a1n a1 vss vss n w=33u l=2.3636u ad='33u*5u+12p' as='33u*5u+12p' pd='33u*2+14u' ps='33u*2+14u'
m7 z sn a0n vss n w=33u l=2.3636u ad='33u*5u+12p' as='33u*5u+12p' pd='33u*2+14u' ps='33u*2+14u'
m8 a1n s z vss n w=33u l=2.3636u ad='33u*5u+12p' as='33u*5u+12p' pd='33u*2+14u' ps='33u*2+14u'
m9 a0n a0 vss vss n w=33u l=2.3636u ad='33u*5u+12p' as='33u*5u+12p' pd='33u*2+14u' ps='33u*2+14u'
m10 sn s vss vss n w=15u l=2.3636u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
.ends
