* Thu Jan 11 12:58:26 CET 2007
.subckt nd2v0x4 a b vdd vss z
*SPICE circuit <nd2v0x4> from XCircuit v3.20

m1 n1 a vss vss n w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m2 z a vdd vdd p w=56u l=2.3636u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m3 z b n1 vss n w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m4 z b vdd vdd p w=56u l=2.3636u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
.ends
