* Spice description of bf1v2x1
* Spice driver version 134999461
* Date 17/05/2007 at  9:05:17
* wsclib 0.13um values
.subckt bf1v2x1 a vdd vss z
M01 an    a     vdd   vdd p  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
M02 an    a     vss   vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M03 vdd   an    z     vdd p  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
M04 vss   an    z     vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
C4  a     vss   0.386f
C1  an    vss   0.430f
C3  z     vss   0.558f
.ends
