* Spice description of iv1_y2
* Spice driver version 134999461
* Date 22/07/2007 at 10:58:37
* vsxlib 0.13um values
.subckt iv1_y2 a vdd vss z
M1  vdd   a     z     vdd p  L=0.12U  W=1.98U  AS=0.5247P   AD=0.5247P   PS=4.49U   PD=4.49U
M2  z     a     vss   vss n  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
C3  a     vss   0.447f
C1  z     vss   0.765f
.ends
