* Thu Jan 11 12:49:16 CET 2007
.subckt iv1v0x8 a vdd vss z
*SPICE circuit <iv1v0x8> from XCircuit v3.20

m1 z a vss vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m2 z a vdd vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
.ends
