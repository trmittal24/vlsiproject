* Fri Apr  8 11:36:53 CEST 2005
.subckt an2v0x6 a b vdd vss z 
*SPICE circuit <an2v0x6> from XCircuit v3.20

m1 z zn vdd vdd p w=81u l=2u ad='81u*5u+12p' as='81u*5u+12p' pd='81u*2+14u' ps='81u*2+14u'
m2 z zn vss vss n w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m3 n1 a vss vss n w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m4 zn a vdd vdd p w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m5 zn b n1 vss n w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m6 zn b vdd vdd p w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
.ends
