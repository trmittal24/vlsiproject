* Tue Aug 10 11:21:07 CEST 2004
.subckt iv1_x1 a vdd vss z 
*SPICE circuit <iv1_x1> from XCircuit v3.10

m1 z a vss vss n w=10u l=2u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m2 z a vdd vdd p w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
.ends
