magic
tech scmos
timestamp 1523182792
<< polysilicon >>
rect 370 -30 372 13
<< metal1 >>
rect -34 228 56 236
rect 270 228 348 233
rect 416 228 447 234
rect 286 195 330 199
rect 417 162 420 164
rect 416 156 420 162
rect 417 155 420 156
rect 631 137 653 143
rect 279 84 283 120
rect 317 88 324 92
rect 279 80 322 84
rect 304 53 308 80
rect 317 42 321 77
rect 285 38 321 42
rect 294 -199 299 38
rect 304 -21 308 21
rect 304 -26 321 -21
rect 304 -192 308 -26
rect 329 -49 333 92
rect 647 73 653 137
rect 527 72 653 73
rect 532 67 653 72
rect 903 33 924 36
rect 438 12 441 26
rect 374 -34 380 -30
rect 304 -196 319 -192
rect 294 -203 321 -199
rect 443 -251 1184 -247
rect -35 -274 59 -265
rect 416 -268 459 -267
rect 272 -273 343 -268
rect 416 -272 458 -268
rect 416 -273 459 -272
<< metal2 >>
rect 280 254 441 259
rect 72 231 76 235
rect 280 195 284 254
rect 362 229 405 233
rect 287 185 324 189
rect 147 77 157 81
rect 208 6 238 10
rect 70 -47 76 -42
rect 287 -69 291 185
rect 287 -78 291 -74
rect 284 -82 291 -78
rect 295 176 323 180
rect 295 -96 299 176
rect 397 156 409 159
rect 362 79 380 83
rect 362 78 376 79
rect 436 72 441 254
rect 886 137 913 141
rect 1148 138 1162 141
rect 436 67 527 72
rect 532 67 533 72
rect 304 25 308 49
rect 629 33 899 36
rect 335 14 339 29
rect 629 29 633 33
rect 441 26 633 29
rect 908 28 913 137
rect 1159 36 1162 138
rect 928 33 1162 36
rect 638 25 913 28
rect 638 21 643 25
rect 311 10 339 14
rect 429 16 643 21
rect 208 -118 220 -113
rect 295 -153 299 -101
rect 282 -157 299 -153
rect 311 -105 315 10
rect 384 5 409 8
rect 429 -21 433 16
rect 320 -26 321 -21
rect 326 -26 433 -21
rect 438 -30 441 8
rect 1257 -8 1268 -4
rect 384 -34 441 -30
rect 353 -47 357 -43
rect 668 -69 669 -67
rect 928 -68 944 -64
rect 928 -69 939 -68
rect 668 -73 672 -69
rect 320 -87 324 -74
rect 928 -77 932 -69
rect 1188 -66 1189 -62
rect 1188 -73 1192 -66
rect 1188 -74 1191 -73
rect 398 -91 424 -87
rect 311 -109 323 -105
rect 154 -199 160 -193
rect 311 -235 315 -109
rect 404 -122 409 -118
rect 364 -147 424 -143
rect 1273 -157 1297 -154
rect 1294 -158 1297 -157
rect 362 -197 376 -193
rect 362 -198 377 -197
rect 373 -201 377 -198
rect 461 -232 462 -231
rect 282 -239 315 -235
rect 399 -251 439 -247
rect 208 -271 239 -268
rect 383 -271 409 -268
rect 458 -268 462 -232
rect 1188 -251 1195 -247
rect 383 -272 412 -271
rect 458 -273 462 -272
<< metal3 >>
rect 75 236 83 237
rect 75 230 76 236
rect 82 230 83 236
rect 75 88 83 230
rect 356 233 363 234
rect 356 229 357 233
rect 362 229 363 233
rect 201 162 209 163
rect 201 156 202 162
rect 208 156 209 162
rect 75 86 147 88
rect 75 84 148 86
rect 75 82 140 84
rect 75 -41 83 82
rect 139 77 140 82
rect 147 77 148 84
rect 139 76 148 77
rect 75 -47 76 -41
rect 82 -47 83 -41
rect 75 -191 83 -47
rect 201 11 209 156
rect 201 6 202 11
rect 208 6 209 11
rect 201 -112 209 6
rect 356 83 363 229
rect 356 78 357 83
rect 362 78 363 83
rect 356 -42 363 78
rect 356 -47 357 -42
rect 362 -47 363 -42
rect 285 -69 326 -68
rect 285 -74 286 -69
rect 291 -74 320 -69
rect 325 -74 326 -69
rect 285 -75 326 -74
rect 335 -95 342 -94
rect 294 -96 336 -95
rect 294 -101 295 -96
rect 300 -100 336 -96
rect 341 -100 342 -95
rect 300 -101 342 -100
rect 294 -102 335 -101
rect 201 -118 202 -112
rect 208 -118 209 -112
rect 75 -193 155 -191
rect 75 -197 147 -193
rect 146 -200 147 -197
rect 154 -200 155 -193
rect 146 -201 155 -200
rect 201 -266 209 -118
rect 356 -193 363 -47
rect 356 -198 357 -193
rect 362 -198 363 -193
rect 356 -199 363 -198
rect 408 159 415 160
rect 408 155 409 159
rect 414 155 415 159
rect 408 9 415 155
rect 408 5 409 9
rect 414 5 415 9
rect 408 -118 415 5
rect 1267 -3 1274 -2
rect 1267 -8 1268 -3
rect 1273 -8 1274 -3
rect 1187 -61 1201 -60
rect 668 -65 680 -64
rect 668 -69 669 -65
rect 674 -69 680 -65
rect 1187 -66 1189 -61
rect 1194 -66 1201 -61
rect 1187 -67 1201 -66
rect 668 -70 680 -69
rect 674 -79 680 -70
rect 938 -68 945 -67
rect 938 -73 939 -68
rect 944 -73 945 -68
rect 938 -74 945 -73
rect 423 -85 680 -79
rect 423 -86 430 -85
rect 423 -91 424 -86
rect 429 -91 430 -86
rect 423 -92 430 -91
rect 939 -103 945 -74
rect 408 -122 409 -118
rect 414 -122 415 -118
rect 201 -272 202 -266
rect 208 -272 209 -266
rect 408 -266 415 -122
rect 423 -110 945 -103
rect 423 -142 430 -110
rect 423 -147 424 -142
rect 429 -147 430 -142
rect 423 -148 430 -147
rect 1194 -247 1201 -67
rect 1267 -152 1274 -8
rect 1267 -157 1268 -152
rect 1273 -157 1274 -152
rect 1267 -158 1274 -157
rect 1194 -251 1195 -247
rect 1200 -251 1201 -247
rect 1194 -252 1201 -251
rect 408 -271 409 -266
rect 414 -271 415 -266
rect 408 -272 415 -271
rect 201 -273 209 -272
<< polycontact >>
rect 370 -34 374 -30
<< m2contact >>
rect 67 231 72 236
rect 405 229 409 233
rect 393 156 397 160
rect 157 77 162 82
rect 304 49 308 53
rect 238 6 242 10
rect 65 -47 70 -42
rect 220 -118 225 -113
rect 160 -199 167 -192
rect 304 21 308 25
rect 321 -26 326 -21
rect 376 75 380 79
rect 527 67 532 72
rect 899 33 903 37
rect 924 33 928 37
rect 437 26 441 30
rect 380 5 384 9
rect 437 8 441 12
rect 380 -34 384 -30
rect 349 -47 353 -43
rect 400 -122 404 -118
rect 1294 -162 1298 -158
rect 377 -201 381 -197
rect 457 -232 461 -228
rect 439 -251 443 -247
rect 1184 -251 1188 -247
rect 239 -271 243 -267
rect 379 -272 383 -268
rect 458 -272 462 -268
<< m3contact >>
rect 76 230 82 236
rect 357 229 362 233
rect 202 156 208 162
rect 140 77 147 84
rect 202 6 208 11
rect 76 -47 82 -41
rect 286 -74 291 -69
rect 409 155 414 159
rect 357 78 362 83
rect 295 -101 300 -96
rect 202 -118 208 -112
rect 409 5 414 9
rect 1268 -8 1273 -3
rect 357 -47 362 -42
rect 669 -69 674 -65
rect 320 -74 325 -69
rect 939 -73 944 -68
rect 1189 -66 1194 -61
rect 424 -91 429 -86
rect 336 -100 341 -95
rect 147 -200 154 -193
rect 409 -122 414 -118
rect 424 -147 429 -142
rect 1268 -157 1273 -152
rect 357 -198 362 -193
rect 202 -272 208 -266
rect 409 -271 414 -266
rect 1195 -251 1200 -247
use decoder  decoder_0
timestamp 1523182792
transform 1 0 58 0 1 160
box -58 -160 229 80
use 3_bitmux  3_bitmux_0
timestamp 1523182792
transform 1 0 347 0 1 159
box -29 -160 85 80
use decoder  decoder_1
timestamp 1523182792
transform 1 0 58 0 1 -117
box -58 -160 229 80
use 3_bitmux  3_bitmux_1
timestamp 1523182792
transform 1 0 347 0 1 -117
box -29 -160 85 80
use subcomp  subcomp_0
timestamp 1523182792
transform 1 0 -477 0 1 40
box 922 -317 2190 330
<< labels >>
rlabel metal1 -32 231 -32 231 3 vdd
rlabel metal1 -30 -270 -30 -270 3 gnd
<< end >>
