* Sat Aug 27 19:28:34 CEST 2005
.subckt nd2v5x8 a b vdd vss z 
*SPICE circuit <nd2v5x8> from XCircuit v3.20

m1 n1 a vss vss n w=72u l=2u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
m2 z a vdd vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
m3 z b n1 vss n w=72u l=2u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
m4 z b vdd vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
.ends
