* Wed Apr  5 08:58:18 CEST 2006
.subckt bf1v0x1 a vdd vss z 
*SPICE circuit <bf1v0x1> from XCircuit v3.20

m1 an a vss vss n w=8u l=2u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
m2 an a vdd vdd p w=13u l=2u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m3 z an vss vss n w=9u l=2u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m4 z an vdd vdd p w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
.ends
