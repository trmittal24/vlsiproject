* Fri Apr  8 11:36:55 CEST 2005
.subckt an2v0x8 a b vdd vss z 
*SPICE circuit <an2v0x8> from XCircuit v3.20

m1 z zn vdd vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
m2 z zn vss vss n w=57u l=2u ad='57u*5u+12p' as='57u*5u+12p' pd='57u*2+14u' ps='57u*2+14u'
m3 n1 a vss vss n w=34u l=2u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
m4 zn a vdd vdd p w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m5 zn b n1 vss n w=34u l=2u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
m6 zn b vdd vdd p w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
.ends
