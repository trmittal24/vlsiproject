* SPICE3 file created from counter.ext - technology: scmos

.include t14y_tsmc_025_level3.txt

M1000 t_0_cp an2v0x3_0_zn t_2_vdd t_2_vdd pfet w=20u l=2u
+ ad=160p pd=56u as=5134p ps=1836u 
M1001 t_2_vdd an2v0x3_0_zn t_0_cp t_2_vdd pfet w=20u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1002 an2v0x3_0_zn an2v0x3_0_a t_2_vdd t_2_vdd pfet w=20u l=2u
+ ad=166p pd=62u as=0p ps=0u 
M1003 t_2_vdd an2v0x3_0_b an2v0x3_0_zn t_2_vdd pfet w=20u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1004 t_2_vss an2v0x3_0_zn t_0_cp t_2_vss nfet w=20u l=2u
+ ad=3631p pd=1406u as=126p ps=54u 
M1005 an2v0x3_0_a_30_9# an2v0x3_0_a t_2_vss t_2_vss nfet w=17u l=2u
+ ad=85p pd=44u as=0p ps=0u 
M1006 an2v0x3_0_zn an2v0x3_0_b an2v0x3_0_a_30_9# t_2_vss nfet w=17u l=2u
+ ad=97p pd=48u as=0p ps=0u 
M1007 t_2_vdd t_0_d t_0_z t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=168p ps=70u 
M1008 t_0_d t_0_n4 t_2_vdd t_2_vdd pfet w=14u l=2u
+ ad=82p pd=42u as=0p ps=0u 
M1009 t_0_a_44_52# t_0_d t_2_vdd t_2_vdd pfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1010 t_0_n4 t_0_ci t_0_a_44_52# t_2_vdd pfet w=6u l=2u
+ ad=78p pd=40u as=0p ps=0u 
M1011 t_0_n2 t_0_cn t_0_n4 t_2_vdd pfet w=12u l=2u
+ ad=96p pd=40u as=0p ps=0u 
M1012 t_2_vdd t_0_n1 t_0_n2 t_2_vdd pfet w=12u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1013 t_0_a_81_58# t_0_n2 t_2_vdd t_2_vdd pfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1014 t_0_n1 t_0_cn t_0_a_81_58# t_2_vdd pfet w=6u l=2u
+ ad=83p pd=42u as=0p ps=0u 
M1015 t_2_vss t_0_d t_0_z t_2_vss nfet w=14u l=2u
+ ad=0p pd=0u as=82p ps=42u 
M1016 t_2_vss t_0_n4 t_0_d t_2_vss nfet w=7u l=2u
+ ad=0p pd=0u as=47p ps=28u 
M1017 t_0_a_98_51# t_0_ci t_0_n1 t_2_vdd pfet w=13u l=2u
+ ad=65p pd=36u as=0p ps=0u 
M1018 t_2_vdd t_0_d t_0_a_98_51# t_2_vdd pfet w=13u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1019 t_0_ci t_0_cn t_2_vdd t_2_vdd pfet w=11u l=2u
+ ad=67p pd=36u as=0p ps=0u 
M1020 t_0_cn t_0_cp t_2_vdd t_2_vdd pfet w=10u l=2u
+ ad=62p pd=34u as=0p ps=0u 
M1021 t_2_vss t_0_cn t_0_ci t_2_vss nfet w=6u l=2u
+ ad=0p pd=0u as=42p ps=26u 
M1022 t_0_a_44_17# t_0_d t_2_vss t_2_vss nfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1023 t_0_n4 t_0_cn t_0_a_44_17# t_2_vss nfet w=6u l=2u
+ ad=48p pd=28u as=0p ps=0u 
M1024 t_0_n2 t_0_ci t_0_n4 t_2_vss nfet w=6u l=2u
+ ad=48p pd=28u as=0p ps=0u 
M1025 t_2_vss t_0_n1 t_0_n2 t_2_vss nfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1026 t_0_a_81_17# t_0_n2 t_2_vss t_2_vss nfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1027 t_0_n1 t_0_ci t_0_a_81_17# t_2_vss nfet w=6u l=2u
+ ad=48p pd=28u as=0p ps=0u 
M1028 t_0_a_98_17# t_0_cn t_0_n1 t_2_vss nfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1029 t_2_vss t_0_d t_0_a_98_17# t_2_vss nfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1030 t_0_cn t_0_cp t_2_vss t_2_vss nfet w=7u l=2u
+ ad=49p pd=28u as=0p ps=0u 
M1031 t_2_vdd bf1v0x6_2_an bf1v0x6_2_z t_2_vdd pfet w=27u l=2u
+ ad=0p pd=0u as=377p ps=138u 
M1032 bf1v0x6_2_z bf1v0x6_2_an t_2_vdd t_2_vdd pfet w=27u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1033 t_2_vdd bf1v0x6_2_an bf1v0x6_2_z t_2_vdd pfet w=27u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1034 bf1v0x6_2_an t_0_z t_2_vdd t_2_vdd pfet w=18u l=2u
+ ad=144p pd=52u as=0p ps=0u 
M1035 t_2_vdd t_0_z bf1v0x6_2_an t_2_vdd pfet w=18u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1036 bf1v0x6_2_z bf1v0x6_2_an t_2_vss t_2_vss nfet w=20u l=2u
+ ad=160p pd=56u as=0p ps=0u 
M1037 t_2_vss bf1v0x6_2_an bf1v0x6_2_z t_2_vss nfet w=20u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1038 bf1v0x6_2_an t_0_z t_2_vss t_2_vss nfet w=19u l=2u
+ ad=121p pd=52u as=0p ps=0u 
M1039 xor2v0x3_0_bn xor2v0x3_1_b t_2_vdd t_2_vdd pfet w=28u l=2u
+ ad=672p pd=216u as=0p ps=0u 
M1040 t_2_vdd xor2v0x3_1_b xor2v0x3_0_bn t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1041 xor2v0x3_0_bn xor2v0x3_1_b t_2_vdd t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1042 t_1_cp xor2v0x3_0_an xor2v0x3_0_bn t_2_vdd pfet w=28u l=2u
+ ad=582p pd=216u as=0p ps=0u 
M1043 xor2v0x3_0_an xor2v0x3_0_bn t_1_cp t_2_vdd pfet w=13u l=2u
+ ad=494p pd=184u as=0p ps=0u 
M1044 t_1_cp xor2v0x3_0_bn xor2v0x3_0_an t_2_vdd pfet w=13u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1045 xor2v0x3_0_bn xor2v0x3_0_an t_1_cp t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1046 t_1_cp xor2v0x3_0_an xor2v0x3_0_bn t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1047 xor2v0x3_0_an xor2v0x3_0_bn t_1_cp t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1048 t_2_vdd t_0_z xor2v0x3_0_an t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1049 xor2v0x3_0_an t_0_z t_2_vdd t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1050 xor2v0x3_0_bn xor2v0x3_1_b t_2_vss t_2_vss nfet w=11u l=2u
+ ad=118p pd=50u as=0p ps=0u 
M1051 t_2_vss xor2v0x3_1_b xor2v0x3_0_bn t_2_vss nfet w=17u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1052 xor2v0x3_0_an xor2v0x3_1_b t_1_cp t_2_vss nfet w=14u l=2u
+ ad=224p pd=88u as=342p ps=148u 
M1053 t_1_cp xor2v0x3_1_b xor2v0x3_0_an t_2_vss nfet w=14u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1054 xor2v0x3_0_a_61_7# xor2v0x3_0_an t_1_cp t_2_vss nfet w=19u l=2u
+ ad=95p pd=48u as=0p ps=0u 
M1055 t_2_vss xor2v0x3_0_bn xor2v0x3_0_a_61_7# t_2_vss nfet w=19u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1056 xor2v0x3_0_a_80_7# xor2v0x3_0_bn t_2_vss t_2_vss nfet w=19u l=2u
+ ad=95p pd=48u as=0p ps=0u 
M1057 t_1_cp xor2v0x3_0_an xor2v0x3_0_a_80_7# t_2_vss nfet w=19u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1058 xor2v0x3_0_an t_0_z t_2_vss t_2_vss nfet w=14u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1059 t_2_vss t_0_z xor2v0x3_0_an t_2_vss nfet w=14u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1060 t_2_vdd t_1_d t_1_z t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=168p ps=70u 
M1061 t_1_d t_1_n4 t_2_vdd t_2_vdd pfet w=14u l=2u
+ ad=82p pd=42u as=0p ps=0u 
M1062 t_1_a_44_52# t_1_d t_2_vdd t_2_vdd pfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1063 t_1_n4 t_1_ci t_1_a_44_52# t_2_vdd pfet w=6u l=2u
+ ad=78p pd=40u as=0p ps=0u 
M1064 t_1_n2 t_1_cn t_1_n4 t_2_vdd pfet w=12u l=2u
+ ad=96p pd=40u as=0p ps=0u 
M1065 t_2_vdd t_1_n1 t_1_n2 t_2_vdd pfet w=12u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1066 t_1_a_81_58# t_1_n2 t_2_vdd t_2_vdd pfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1067 t_1_n1 t_1_cn t_1_a_81_58# t_2_vdd pfet w=6u l=2u
+ ad=83p pd=42u as=0p ps=0u 
M1068 t_2_vss t_1_d t_1_z t_2_vss nfet w=14u l=2u
+ ad=0p pd=0u as=82p ps=42u 
M1069 t_2_vss t_1_n4 t_1_d t_2_vss nfet w=7u l=2u
+ ad=0p pd=0u as=47p ps=28u 
M1070 t_1_a_98_51# t_1_ci t_1_n1 t_2_vdd pfet w=13u l=2u
+ ad=65p pd=36u as=0p ps=0u 
M1071 t_2_vdd t_1_d t_1_a_98_51# t_2_vdd pfet w=13u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1072 t_1_ci t_1_cn t_2_vdd t_2_vdd pfet w=11u l=2u
+ ad=67p pd=36u as=0p ps=0u 
M1073 t_1_cn t_1_cp t_2_vdd t_2_vdd pfet w=10u l=2u
+ ad=62p pd=34u as=0p ps=0u 
M1074 t_2_vss t_1_cn t_1_ci t_2_vss nfet w=6u l=2u
+ ad=0p pd=0u as=42p ps=26u 
M1075 t_1_a_44_17# t_1_d t_2_vss t_2_vss nfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1076 t_1_n4 t_1_cn t_1_a_44_17# t_2_vss nfet w=6u l=2u
+ ad=48p pd=28u as=0p ps=0u 
M1077 t_1_n2 t_1_ci t_1_n4 t_2_vss nfet w=6u l=2u
+ ad=48p pd=28u as=0p ps=0u 
M1078 t_2_vss t_1_n1 t_1_n2 t_2_vss nfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1079 t_1_a_81_17# t_1_n2 t_2_vss t_2_vss nfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1080 t_1_n1 t_1_ci t_1_a_81_17# t_2_vss nfet w=6u l=2u
+ ad=48p pd=28u as=0p ps=0u 
M1081 t_1_a_98_17# t_1_cn t_1_n1 t_2_vss nfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1082 t_2_vss t_1_d t_1_a_98_17# t_2_vss nfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1083 t_1_cn t_1_cp t_2_vss t_2_vss nfet w=7u l=2u
+ ad=49p pd=28u as=0p ps=0u 
M1084 t_2_vdd bf1v0x6_1_an bf1v0x6_1_z t_2_vdd pfet w=27u l=2u
+ ad=0p pd=0u as=377p ps=138u 
M1085 bf1v0x6_1_z bf1v0x6_1_an t_2_vdd t_2_vdd pfet w=27u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1086 t_2_vdd bf1v0x6_1_an bf1v0x6_1_z t_2_vdd pfet w=27u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1087 bf1v0x6_1_an t_1_z t_2_vdd t_2_vdd pfet w=18u l=2u
+ ad=144p pd=52u as=0p ps=0u 
M1088 t_2_vdd t_1_z bf1v0x6_1_an t_2_vdd pfet w=18u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1089 bf1v0x6_1_z bf1v0x6_1_an t_2_vss t_2_vss nfet w=20u l=2u
+ ad=160p pd=56u as=0p ps=0u 
M1090 t_2_vss bf1v0x6_1_an bf1v0x6_1_z t_2_vss nfet w=20u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1091 bf1v0x6_1_an t_1_z t_2_vss t_2_vss nfet w=19u l=2u
+ ad=121p pd=52u as=0p ps=0u 
M1092 xor2v0x3_1_bn xor2v0x3_1_b t_2_vdd t_2_vdd pfet w=28u l=2u
+ ad=672p pd=216u as=0p ps=0u 
M1093 t_2_vdd xor2v0x3_1_b xor2v0x3_1_bn t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1094 xor2v0x3_1_bn xor2v0x3_1_b t_2_vdd t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1095 t_2_cp xor2v0x3_1_an xor2v0x3_1_bn t_2_vdd pfet w=28u l=2u
+ ad=582p pd=216u as=0p ps=0u 
M1096 xor2v0x3_1_an xor2v0x3_1_bn t_2_cp t_2_vdd pfet w=13u l=2u
+ ad=494p pd=184u as=0p ps=0u 
M1097 t_2_cp xor2v0x3_1_bn xor2v0x3_1_an t_2_vdd pfet w=13u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1098 xor2v0x3_1_bn xor2v0x3_1_an t_2_cp t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1099 t_2_cp xor2v0x3_1_an xor2v0x3_1_bn t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1100 xor2v0x3_1_an xor2v0x3_1_bn t_2_cp t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1101 t_2_vdd t_1_z xor2v0x3_1_an t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1102 xor2v0x3_1_an t_1_z t_2_vdd t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1103 xor2v0x3_1_bn xor2v0x3_1_b t_2_vss t_2_vss nfet w=11u l=2u
+ ad=118p pd=50u as=0p ps=0u 
M1104 t_2_vss xor2v0x3_1_b xor2v0x3_1_bn t_2_vss nfet w=17u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1105 xor2v0x3_1_an xor2v0x3_1_b t_2_cp t_2_vss nfet w=14u l=2u
+ ad=224p pd=88u as=342p ps=148u 
M1106 t_2_cp xor2v0x3_1_b xor2v0x3_1_an t_2_vss nfet w=14u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1107 xor2v0x3_1_a_61_7# xor2v0x3_1_an t_2_cp t_2_vss nfet w=19u l=2u
+ ad=95p pd=48u as=0p ps=0u 
M1108 t_2_vss xor2v0x3_1_bn xor2v0x3_1_a_61_7# t_2_vss nfet w=19u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1109 xor2v0x3_1_a_80_7# xor2v0x3_1_bn t_2_vss t_2_vss nfet w=19u l=2u
+ ad=95p pd=48u as=0p ps=0u 
M1110 t_2_cp xor2v0x3_1_an xor2v0x3_1_a_80_7# t_2_vss nfet w=19u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1111 xor2v0x3_1_an t_1_z t_2_vss t_2_vss nfet w=14u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1112 t_2_vss t_1_z xor2v0x3_1_an t_2_vss nfet w=14u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1113 t_2_vdd t_2_d t_2_z t_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=168p ps=70u 
M1114 t_2_d t_2_n4 t_2_vdd t_2_vdd pfet w=14u l=2u
+ ad=82p pd=42u as=0p ps=0u 
M1115 t_2_a_44_52# t_2_d t_2_vdd t_2_vdd pfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1116 t_2_n4 t_2_ci t_2_a_44_52# t_2_vdd pfet w=6u l=2u
+ ad=78p pd=40u as=0p ps=0u 
M1117 t_2_n2 t_2_cn t_2_n4 t_2_vdd pfet w=12u l=2u
+ ad=96p pd=40u as=0p ps=0u 
M1118 t_2_vdd t_2_n1 t_2_n2 t_2_vdd pfet w=12u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1119 t_2_a_81_58# t_2_n2 t_2_vdd t_2_vdd pfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1120 t_2_n1 t_2_cn t_2_a_81_58# t_2_vdd pfet w=6u l=2u
+ ad=83p pd=42u as=0p ps=0u 
M1121 t_2_vss t_2_d t_2_z t_2_vss nfet w=14u l=2u
+ ad=0p pd=0u as=82p ps=42u 
M1122 t_2_vss t_2_n4 t_2_d t_2_vss nfet w=7u l=2u
+ ad=0p pd=0u as=47p ps=28u 
M1123 t_2_a_98_51# t_2_ci t_2_n1 t_2_vdd pfet w=13u l=2u
+ ad=65p pd=36u as=0p ps=0u 
M1124 t_2_vdd t_2_d t_2_a_98_51# t_2_vdd pfet w=13u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1125 t_2_ci t_2_cn t_2_vdd t_2_vdd pfet w=11u l=2u
+ ad=67p pd=36u as=0p ps=0u 
M1126 t_2_cn t_2_cp t_2_vdd t_2_vdd pfet w=10u l=2u
+ ad=62p pd=34u as=0p ps=0u 
M1127 t_2_vss t_2_cn t_2_ci t_2_vss nfet w=6u l=2u
+ ad=0p pd=0u as=42p ps=26u 
M1128 t_2_a_44_17# t_2_d t_2_vss t_2_vss nfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1129 t_2_n4 t_2_cn t_2_a_44_17# t_2_vss nfet w=6u l=2u
+ ad=48p pd=28u as=0p ps=0u 
M1130 t_2_n2 t_2_ci t_2_n4 t_2_vss nfet w=6u l=2u
+ ad=48p pd=28u as=0p ps=0u 
M1131 t_2_vss t_2_n1 t_2_n2 t_2_vss nfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1132 t_2_a_81_17# t_2_n2 t_2_vss t_2_vss nfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1133 t_2_n1 t_2_ci t_2_a_81_17# t_2_vss nfet w=6u l=2u
+ ad=48p pd=28u as=0p ps=0u 
M1134 t_2_a_98_17# t_2_cn t_2_n1 t_2_vss nfet w=6u l=2u
+ ad=30p pd=22u as=0p ps=0u 
M1135 t_2_vss t_2_d t_2_a_98_17# t_2_vss nfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1136 t_2_cn t_2_cp t_2_vss t_2_vss nfet w=7u l=2u
+ ad=49p pd=28u as=0p ps=0u 
M1137 t_2_vdd bf1v0x6_0_an bf1v0x6_0_z t_2_vdd pfet w=27u l=2u
+ ad=0p pd=0u as=377p ps=138u 
M1138 bf1v0x6_0_z bf1v0x6_0_an t_2_vdd t_2_vdd pfet w=27u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1139 t_2_vdd bf1v0x6_0_an bf1v0x6_0_z t_2_vdd pfet w=27u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1140 bf1v0x6_0_an t_2_z t_2_vdd t_2_vdd pfet w=18u l=2u
+ ad=144p pd=52u as=0p ps=0u 
M1141 t_2_vdd t_2_z bf1v0x6_0_an t_2_vdd pfet w=18u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1142 bf1v0x6_0_z bf1v0x6_0_an t_2_vss t_2_vss nfet w=20u l=2u
+ ad=160p pd=56u as=0p ps=0u 
M1143 t_2_vss bf1v0x6_0_an bf1v0x6_0_z t_2_vss nfet w=20u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1144 bf1v0x6_0_an t_2_z t_2_vss t_2_vss nfet w=19u l=2u
+ ad=121p pd=52u as=0p ps=0u 
C0 t_2_vdd t_1_z 28.2fF
C1 t_2_vdd bf1v0x6_2_an 15.4fF
C2 t_2_vss t_0_z 21.0fF
C3 xor2v0x3_0_bn t_1_cp 7.1fF
C4 an2v0x3_0_b t_2_vss 5.5fF
C5 t_2_n2 t_2_vdd 12.4fF
C6 t_0_ci t_2_vdd 16.6fF
C7 xor2v0x3_1_b t_2_vss 51.1fF
C8 t_0_cn t_2_vss 17.1fF
C9 t_2_vss bf1v0x6_0_an 11.0fF
C10 t_2_vss t_1_ci 27.5fF
C11 t_2_vdd t_2_z 17.5fF
C12 an2v0x3_0_a t_2_vss 6.3fF
C13 t_0_n4 t_2_vss 7.3fF
C14 t_2_vdd t_0_z 28.1fF
C15 t_2_vss bf1v0x6_1_z 3.5fF
C16 xor2v0x3_1_an t_2_cp 3.6fF
C17 an2v0x3_0_b t_2_vdd 6.5fF
C18 xor2v0x3_0_an t_1_cp 3.6fF
C19 xor2v0x3_1_b t_2_vdd 38.6fF
C20 t_0_cn t_2_vdd 46.5fF
C21 t_2_vdd bf1v0x6_0_an 15.4fF
C22 t_2_vdd t_1_ci 16.6fF
C23 t_2_vss t_2_n4 7.3fF
C24 xor2v0x3_0_bn t_2_vss 12.6fF
C25 xor2v0x3_1_an t_2_vss 18.3fF
C26 an2v0x3_0_a t_2_vdd 5.3fF
C27 t_2_vss t_1_n2 7.2fF
C28 t_2_cn t_2_vss 17.1fF
C29 t_0_n4 t_2_vdd 8.9fF
C30 t_2_vdd bf1v0x6_1_z 3.9fF
C31 t_2_ci t_2_vss 27.5fF
C32 t_2_vss bf1v0x6_0_z 3.5fF
C33 t_2_vdd t_2_n4 8.9fF
C34 t_2_vdd xor2v0x3_0_bn 24.1fF
C35 xor2v0x3_1_an t_2_vdd 19.1fF
C36 t_2_d t_2_vss 28.2fF
C37 xor2v0x3_0_an t_2_vss 18.3fF
C38 t_2_vdd t_1_n2 12.4fF
C39 t_2_cn t_2_vdd 46.5fF
C40 t_2_vss t_1_n1 9.9fF
C41 t_2_vss bf1v0x6_2_z 3.5fF
C42 bf1v0x6_1_an t_2_vss 11.0fF
C43 t_2_vdd t_2_ci 16.6fF
C44 t_2_vdd bf1v0x6_0_z 3.9fF
C45 t_0_cp t_2_vss 4.7fF
C46 t_0_n1 t_2_vss 9.9fF
C47 t_2_vdd t_2_d 18.0fF
C48 xor2v0x3_0_an t_2_vdd 19.1fF
C49 t_2_vss t_0_n2 7.2fF
C50 t_2_vss t_1_cp 9.0fF
C51 t_2_vdd t_1_n1 8.4fF
C52 t_2_vdd bf1v0x6_2_z 3.9fF
C53 t_2_n1 t_2_vss 9.9fF
C54 t_2_vss an2v0x3_0_zn 9.5fF
C55 t_2_vdd bf1v0x6_1_an 15.4fF
C56 t_0_d t_2_vss 28.2fF
C57 t_0_cp t_2_vdd 18.8fF
C58 xor2v0x3_1_bn t_2_cp 8.8fF
C59 t_2_vss t_1_n4 7.3fF
C60 t_2_vdd t_0_n1 8.4fF
C61 t_0_d t_0_ci 4.2fF
C62 t_1_d t_2_vss 28.2fF
C63 t_1_cn t_2_vss 17.1fF
C64 t_2_vdd t_0_n2 12.4fF
C65 t_2_cp t_2_vss 9.0fF
C66 t_2_vdd t_1_cp 22.3fF
C67 xor2v0x3_1_bn t_2_vss 12.6fF
C68 t_2_vss t_1_z 20.7fF
C69 t_2_vss bf1v0x6_2_an 11.0fF
C70 t_2_n1 t_2_vdd 8.4fF
C71 t_2_vdd an2v0x3_0_zn 13.3fF
C72 t_0_d t_2_vdd 18.0fF
C73 t_2_n2 t_2_vss 7.2fF
C74 t_2_vdd t_1_n4 8.9fF
C75 t_0_ci t_2_vss 27.5fF
C76 t_1_d t_2_vdd 18.0fF
C77 t_2_vdd t_1_cn 46.5fF
C78 t_2_cp t_2_vdd 23.0fF
C79 t_2_vss t_2_z 10.3fF
C80 t_1_d t_1_ci 4.2fF
C81 t_2_d t_2_ci 4.2fF
C82 xor2v0x3_1_b t_2_cp 6.8fF
C83 xor2v0x3_1_bn t_2_vdd 24.1fF
C84 t_2_vss 0 335.3fF
C85 t_2_vdd 0 40.8fF


v_dd t_2_vdd 0 5
v_ss t_2_vss 0 0
v_gg_cp an2v0x3_0_a 0 PULSE(0 5 0 0.1n 0.1n 30n 60n)
v_dd_en an2v0x3_0_b 0 PULSE(5 0 200n 0.1n 0.1n 200n 400n)
v_dd_ud xor2v0x3_1_b 0 0

.control
 tran 1n 800n
 plot (an2v0x3_0_a + 5) (t_0_z) (bf1v0x6_2_z - 5) (bf1v0x6_1_z - 10) ( bf1v0x6_0_z - 15) (an2v0x3_0_b - 20)
.endc

.end