* Tue Aug 10 11:21:07 CEST 2004
.subckt cgn2_x4 a b c vdd vss z 
*SPICE circuit <cgn2_x4> from XCircuit v3.10

m1 z zn vss vss n w=37u l=2u ad='37u*5u+12p' as='37u*5u+12p' pd='37u*2+14u' ps='37u*2+14u'
m2 zn b n4 vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m3 z zn vdd vdd p w=74u l=2u ad='74u*5u+12p' as='74u*5u+12p' pd='74u*2+14u' ps='74u*2+14u'
m4 n4 a vss vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m5 n3 b vss vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m6 zn c n3 vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m7 zn b n2 vdd p w=62u l=2u ad='62u*5u+12p' as='62u*5u+12p' pd='62u*2+14u' ps='62u*2+14u'
m8 n2 a vdd vdd p w=62u l=2u ad='62u*5u+12p' as='62u*5u+12p' pd='62u*2+14u' ps='62u*2+14u'
m9 zn c n1 vdd p w=62u l=2u ad='62u*5u+12p' as='62u*5u+12p' pd='62u*2+14u' ps='62u*2+14u'
m10 n1 b vdd vdd p w=62u l=2u ad='62u*5u+12p' as='62u*5u+12p' pd='62u*2+14u' ps='62u*2+14u'
m11 n1 a vdd vdd p w=62u l=2u ad='62u*5u+12p' as='62u*5u+12p' pd='62u*2+14u' ps='62u*2+14u'
m12 n3 a vss vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
.ends
