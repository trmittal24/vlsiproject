* Mon Aug 16 14:22:56 CEST 2004
.subckt buf_x8 i q vdd vss 
*SPICE circuit <buf_x8> from XCircuit v3.10

m1 in i vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m2 in i vdd vdd p w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m3 q in vss vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m4 q in vdd vdd p w=160u l=2u ad='160u*5u+12p' as='160u*5u+12p' pd='160u*2+14u' ps='160u*2+14u'
.ends
