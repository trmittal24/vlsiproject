* Tue Aug 10 11:21:07 CEST 2004
.subckt oan21_x1 a1 a2 b vdd vss z 
*SPICE circuit <oan21_x1> from XCircuit v3.10

m1 z zn vss vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m2 z zn vdd vdd p w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m3 n1 a1 vdd vdd p w=26u l=2.3636u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m4 zn b vdd vdd p w=14u l=2.3636u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m5 ext16 a2 ext17 vss n w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m6 n2 b vss vss n w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m7 zn a1 n2 vss n w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m8 zn a2 n1 vdd p w=26u l=2.3636u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
.ends
