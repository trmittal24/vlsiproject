* Spice description of bf1v0x2
* Spice driver version 134999461
* Date 17/05/2007 at  9:04:29
* vsclib 0.13um values
.subckt bf1v0x2 a vdd vss z
M01 an    a     vdd   vdd p  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
M02 an    a     vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
M03 vdd   an    z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M04 vss   an    z     vss n  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
C4  a     vss   0.321f
C3  an    vss   0.460f
C2  z     vss   1.111f
.ends
