* Tue Aug 10 11:21:07 CEST 2004
.subckt iv1_x3 a vdd vss z 
*SPICE circuit <iv1_x3> from XCircuit v3.10

m1 z a vss vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m2 z a vdd vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
.ends
