* Mon Aug 16 14:10:59 CEST 2004
.subckt nd2v0x6 a b vdd vss z 
*SPICE circuit <nd2v0x6> from XCircuit v3.10

m1 n1 a vss vss n w=60u l=2u ad='60u*5u+12p' as='60u*5u+12p' pd='60u*2+14u' ps='60u*2+14u'
m2 z a vdd vdd p w=72u l=2u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
m3 z b n1 vss n w=60u l=2u ad='60u*5u+12p' as='60u*5u+12p' pd='60u*2+14u' ps='60u*2+14u'
m4 z b vdd vdd p w=72u l=2u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
.ends
