* Fri Apr  7 16:04:48 CEST 2006
.subckt aoi21v0x05 a1 a2 b vdd vss z 
*SPICE circuit <aoi21v0x05> from XCircuit v3.20

m1 n1 a2 vdd vdd p w=17u l=2u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m2 n1 a1 vdd vdd p w=17u l=2u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m3 n2 a1 vss vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m4 z b vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m5 z a2 n2 vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m6 z b n1 vdd p w=17u l=2u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
.ends
