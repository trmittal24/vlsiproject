* Spice description of nr2v1x05
* Spice driver version 134999461
* Date 17/05/2007 at  9:26:26
* vsclib 0.13um values
.subckt nr2v1x05 a b vdd vss z
M01 vdd   a     n1    vdd p  L=0.12U  W=0.825U AS=0.218625P AD=0.218625P PS=2.18U   PD=2.18U
M02 vss   a     z     vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M03 n1    b     z     vdd p  L=0.12U  W=0.825U AS=0.218625P AD=0.218625P PS=2.18U   PD=2.18U
M04 z     b     vss   vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
C4  a     vss   0.379f
C3  b     vss   0.330f
C1  z     vss   0.616f
.ends
