* Mon Aug 16 14:10:58 CEST 2004
.subckt iv1v1x1 a vdd vss z 
*SPICE circuit <iv1v1x1> from XCircuit v3.10

m1 z a vss vss n w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m2 z a vdd vdd p w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
.ends
