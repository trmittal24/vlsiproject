* Spice description of nr3_x05
* Spice driver version 134999461
* Date 22/07/2007 at 10:59:31
* vsxlib 0.13um values
.subckt nr3_x05 a b c vdd vss z
M1  n2    c     z     vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M2  n1    b     n2    vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M3  vdd   a     n1    vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M4  z     c     vss   vss n  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M5  vss   b     z     vss n  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M6  z     a     vss   vss n  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
C5  a     vss   0.553f
C3  b     vss   0.620f
C4  c     vss   0.702f
C2  z     vss   0.862f
.ends
