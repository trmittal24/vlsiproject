* Spice description of o3_x2
* Spice driver version 134999461
* Date 21/07/2007 at 19:31:33
* sxlib 0.13um values
.subckt o3_x2 i0 i1 i2 q vdd vss
Mtr_00001 sig3  i2    vss   vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00002 sig3  i0    vss   vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00003 vss   i1    sig3  vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00004 vss   sig3  q     vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00005 vdd   i0    sig5  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00006 sig5  i1    sig6  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00007 sig6  i2    sig3  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00008 q     sig3  vdd   vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
C8  i0    vss   0.668f
C7  i1    vss   0.668f
C9  i2    vss   0.645f
C1  q     vss   1.066f
C3  sig3  vss   1.049f
.ends
