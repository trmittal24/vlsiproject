* Spice description of iv1_x4
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:10
*
.subckt iv1_x4 a vdd vss z 
M1  z     a     vdd   vdd p  L=0.13U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U  
M2  vdd   a     z     vdd p  L=0.13U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U  
M3  vss   a     z     vss n  L=0.13U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U  
M4  z     a     vss   vss n  L=0.13U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U  
C4  a     vss   1.313f
C3  vdd   vss   1.468f
C1  z     vss   2.641f
.ends
