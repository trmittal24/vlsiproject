* Spice description of nd2v0x2
* Spice driver version 134999461
* Date 17/06/2007 at 14:03:11
* vgalib 0.13um values
.subckt nd2v0x2 a b vdd vss z
Mtr_00001 sig1  a     vss   vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00002 z     b     sig1  vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00003 vdd   b     z     vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
Mtr_00004 z     a     vdd   vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
C4  a     vss   0.508f
C5  b     vss   0.535f
C2  z     vss   0.921f
.ends
