* Tue Feb 20 08:57:11 CET 2007
.subckt iv1v6x2 a vdd vss z
*SPICE circuit <iv1v6x2> from XCircuit v3.20

m1 z a vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m2 z a vdd vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
.ends
