* Sat Apr  9 11:13:27 CEST 2005
.subckt nr2av0x3 a b vdd vss z 
*SPICE circuit <nr2av0x3> from XCircuit v3.20

m1 an a vss vss n w=14u l=2u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m2 an a vdd vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m3 z an vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m4 n1 an vdd vdd p w=75u l=2u ad='75u*5u+12p' as='75u*5u+12p' pd='75u*2+14u' ps='75u*2+14u'
m5 z b vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m6 z b n1 vdd p w=75u l=2u ad='75u*5u+12p' as='75u*5u+12p' pd='75u*2+14u' ps='75u*2+14u'
.ends
