* Spice description of aoi21bv0x05
* Spice driver version 134999461
* Date 17/05/2007 at  9:00:51
* wsclib 0.13um values
.subckt aoi21bv0x05 a1 a2 b vdd vss z
M01 n1    a1    vdd   vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M02 vss   a1    n2    vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M03 vdd   a2    n1    vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M04 n2    a2    z     vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M05 n1    06    z     vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M06 z     06    vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M07 vdd   b     06    vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M08 06    b     vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
C5  06    vss   0.579f
C6  a1    vss   0.460f
C4  a2    vss   0.441f
C7  b     vss   0.577f
C9  n1    vss   0.220f
C2  z     vss   0.698f
.ends
