* Mon Aug 16 14:10:58 CEST 2004
.subckt iv1v0x3 a vdd vss z 
*SPICE circuit <iv1v0x3> from XCircuit v3.10

m1 z a vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m2 z a vdd vdd p w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
.ends
