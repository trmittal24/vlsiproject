* SPICE3 file created from comp.ext - technology: scmos

.include t14y_tsmc_025_level3.txt

M1000 nd3v0x2_0_z nr3v0x2_0_z an3v0x2_2_vdd an3v0x2_2_w_n4_32# pfet w=14u l=2u
+ ad=392p pd=120u as=7344p ps=2472u 
M1001 an3v0x2_2_vdd nr3v0x2_0_z nd3v0x2_0_z an3v0x2_2_w_n4_32# pfet w=14u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1002 nd3v0x2_0_z nd3v0x2_0_c an3v0x2_2_vdd an3v0x2_2_w_n4_32# pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1003 an3v0x2_2_vdd nd3v0x2_0_a nd3v0x2_0_z an3v0x2_2_w_n4_32# pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1004 nd3v0x2_0_a_14_12# nd3v0x2_0_a an2v0x2_0_vss an2v0x2_0_vss nfet w=14u l=2u
+ ad=70p pd=38u as=4084p ps=1438u 
M1005 nd3v0x2_0_a_21_12# nr3v0x2_0_z nd3v0x2_0_a_14_12# an2v0x2_0_vss nfet w=14u l=2u
+ ad=70p pd=38u as=0p ps=0u 
M1006 nd3v0x2_0_z nd3v0x2_0_c nd3v0x2_0_a_21_12# an2v0x2_0_vss nfet w=14u l=2u
+ ad=112p pd=44u as=0p ps=0u 
M1007 nd3v0x2_0_a_38_12# nd3v0x2_0_c nd3v0x2_0_z an2v0x2_0_vss nfet w=14u l=2u
+ ad=70p pd=38u as=0p ps=0u 
M1008 nd3v0x2_0_a_45_12# nr3v0x2_0_z nd3v0x2_0_a_38_12# an2v0x2_0_vss nfet w=14u l=2u
+ ad=70p pd=38u as=0p ps=0u 
M1009 an2v0x2_0_vss nd3v0x2_0_a nd3v0x2_0_a_45_12# an2v0x2_0_vss nfet w=14u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1010 an3v0x2_2_vdd an3v0x2_1_zn nr2v0x2_1_a an3v0x2_2_w_n4_32# pfet w=28u l=2u
+ ad=0p pd=0u as=166p ps=70u 
M1011 an3v0x2_1_zn an3v0x2_1_a an3v0x2_2_vdd an3v0x2_2_w_n4_32# pfet w=17u l=2u
+ ad=233p pd=98u as=0p ps=0u 
M1012 an3v0x2_2_vdd an3v0x2_2_b an3v0x2_1_zn an3v0x2_2_w_n4_32# pfet w=17u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1013 an3v0x2_1_zn an3v0x2_2_c an3v0x2_2_vdd an3v0x2_2_w_n4_32# pfet w=17u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1014 an2v0x2_0_vss an3v0x2_1_zn nr2v0x2_1_a an2v0x2_0_vss nfet w=14u l=2u
+ ad=0p pd=0u as=82p ps=42u 
M1015 an3v0x2_1_a_24_8# an3v0x2_1_a an2v0x2_0_vss an2v0x2_0_vss nfet w=17u l=2u
+ ad=85p pd=44u as=0p ps=0u 
M1016 an3v0x2_1_a_31_8# an3v0x2_2_b an3v0x2_1_a_24_8# an2v0x2_0_vss nfet w=17u l=2u
+ ad=85p pd=44u as=0p ps=0u 
M1017 an3v0x2_1_zn an3v0x2_2_c an3v0x2_1_a_31_8# an2v0x2_0_vss nfet w=17u l=2u
+ ad=97p pd=48u as=0p ps=0u 
M1018 nr3v0x2_0_a_13_39# an3v0x2_2_z nr3v0x2_0_z an3v0x2_2_w_n4_32# pfet w=27u l=2u
+ ad=135p pd=64u as=377p ps=138u 
M1019 nr3v0x2_0_a_20_39# an3v0x2_0_z nr3v0x2_0_a_13_39# an3v0x2_2_w_n4_32# pfet w=27u l=2u
+ ad=135p pd=64u as=0p ps=0u 
M1020 an3v0x2_2_vdd nr3v0x2_0_a nr3v0x2_0_a_20_39# an3v0x2_2_w_n4_32# pfet w=27u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1021 nr3v0x2_0_a_37_39# nr3v0x2_0_a an3v0x2_2_vdd an3v0x2_2_w_n4_32# pfet w=27u l=2u
+ ad=135p pd=64u as=0p ps=0u 
M1022 nr3v0x2_0_a_44_39# an3v0x2_0_z nr3v0x2_0_a_37_39# an3v0x2_2_w_n4_32# pfet w=27u l=2u
+ ad=135p pd=64u as=0p ps=0u 
M1023 nr3v0x2_0_z an3v0x2_2_z nr3v0x2_0_a_44_39# an3v0x2_2_w_n4_32# pfet w=27u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1024 nr3v0x2_0_a_61_39# an3v0x2_2_z nr3v0x2_0_z an3v0x2_2_w_n4_32# pfet w=27u l=2u
+ ad=135p pd=64u as=0p ps=0u 
M1025 nr3v0x2_0_a_68_39# an3v0x2_0_z nr3v0x2_0_a_61_39# an3v0x2_2_w_n4_32# pfet w=27u l=2u
+ ad=135p pd=64u as=0p ps=0u 
M1026 an3v0x2_2_vdd nr3v0x2_0_a nr3v0x2_0_a_68_39# an3v0x2_2_w_n4_32# pfet w=27u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1027 an2v0x2_0_vss an3v0x2_2_z nr3v0x2_0_z an2v0x2_0_vss nfet w=15u l=2u
+ ad=0p pd=0u as=207p ps=90u 
M1028 nr3v0x2_0_z an3v0x2_0_z an2v0x2_0_vss an2v0x2_0_vss nfet w=15u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1029 an2v0x2_0_vss nr3v0x2_0_a nr3v0x2_0_z an2v0x2_0_vss nfet w=15u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1030 an3v0x2_2_vdd an3v0x2_2_zn an3v0x2_2_z an3v0x2_2_w_n4_32# pfet w=28u l=2u
+ ad=0p pd=0u as=166p ps=70u 
M1031 an3v0x2_2_zn an3v0x2_2_a an3v0x2_2_vdd an3v0x2_2_w_n4_32# pfet w=17u l=2u
+ ad=233p pd=98u as=0p ps=0u 
M1032 an3v0x2_2_vdd an3v0x2_2_b an3v0x2_2_zn an3v0x2_2_w_n4_32# pfet w=17u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1033 an3v0x2_2_zn an3v0x2_2_c an3v0x2_2_vdd an3v0x2_2_w_n4_32# pfet w=17u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1034 an2v0x2_0_vss an3v0x2_2_zn an3v0x2_2_z an2v0x2_0_vss nfet w=14u l=2u
+ ad=0p pd=0u as=82p ps=42u 
M1035 an3v0x2_2_a_24_8# an3v0x2_2_a an2v0x2_0_vss an2v0x2_0_vss nfet w=17u l=2u
+ ad=85p pd=44u as=0p ps=0u 
M1036 an3v0x2_2_a_31_8# an3v0x2_2_b an3v0x2_2_a_24_8# an2v0x2_0_vss nfet w=17u l=2u
+ ad=85p pd=44u as=0p ps=0u 
M1037 an3v0x2_2_zn an3v0x2_2_c an3v0x2_2_a_31_8# an2v0x2_0_vss nfet w=17u l=2u
+ ad=97p pd=48u as=0p ps=0u 
M1038 nr2v0x2_1_a_11_39# nr2v0x2_1_a an3v0x2_2_vdd an3v0x2_2_vdd pfet w=27u l=2u
+ ad=135p pd=64u as=0p ps=0u 
M1039 nd3v0x2_0_c an3v0x2_3_z nr2v0x2_1_a_11_39# an3v0x2_2_vdd pfet w=27u l=2u
+ ad=216p pd=70u as=0p ps=0u 
M1040 nr2v0x2_1_a_28_39# an3v0x2_3_z nd3v0x2_0_c an3v0x2_2_vdd pfet w=27u l=2u
+ ad=135p pd=64u as=0p ps=0u 
M1041 an3v0x2_2_vdd nr2v0x2_1_a nr2v0x2_1_a_28_39# an3v0x2_2_vdd pfet w=27u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1042 nd3v0x2_0_c nr2v0x2_1_a an2v0x2_0_vss an2v0x2_0_vss nfet w=15u l=2u
+ ad=120p pd=46u as=0p ps=0u 
M1043 an2v0x2_0_vss an3v0x2_3_z nd3v0x2_0_c an2v0x2_0_vss nfet w=15u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1044 an3v0x2_2_vdd an3v0x2_3_zn an3v0x2_3_z an3v0x2_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=166p ps=70u 
M1045 an3v0x2_3_zn an2v0x2_0_b an3v0x2_2_vdd an3v0x2_2_vdd pfet w=17u l=2u
+ ad=233p pd=98u as=0p ps=0u 
M1046 an3v0x2_2_vdd an3v0x2_0_b an3v0x2_3_zn an3v0x2_2_vdd pfet w=17u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1047 an3v0x2_3_zn an3v0x2_2_a an3v0x2_2_vdd an3v0x2_2_vdd pfet w=17u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1048 an2v0x2_0_vss an3v0x2_3_zn an3v0x2_3_z an2v0x2_0_vss nfet w=14u l=2u
+ ad=0p pd=0u as=82p ps=42u 
M1049 an3v0x2_3_a_24_8# an2v0x2_0_b an2v0x2_0_vss an2v0x2_0_vss nfet w=17u l=2u
+ ad=85p pd=44u as=0p ps=0u 
M1050 an3v0x2_3_a_31_8# an3v0x2_0_b an3v0x2_3_a_24_8# an2v0x2_0_vss nfet w=17u l=2u
+ ad=85p pd=44u as=0p ps=0u 
M1051 an3v0x2_3_zn an3v0x2_2_a an3v0x2_3_a_31_8# an2v0x2_0_vss nfet w=17u l=2u
+ ad=97p pd=48u as=0p ps=0u 
M1052 an3v0x2_2_vdd an3v0x2_0_zn an3v0x2_0_z an3v0x2_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=166p ps=70u 
M1053 an3v0x2_0_zn an3v0x2_1_a an3v0x2_2_vdd an3v0x2_2_vdd pfet w=17u l=2u
+ ad=233p pd=98u as=0p ps=0u 
M1054 an3v0x2_2_vdd an3v0x2_0_b an3v0x2_0_zn an3v0x2_2_vdd pfet w=17u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1055 an3v0x2_0_zn an2v0x2_0_b an3v0x2_2_vdd an3v0x2_2_vdd pfet w=17u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1056 an2v0x2_0_vss an3v0x2_0_zn an3v0x2_0_z an2v0x2_0_vss nfet w=14u l=2u
+ ad=0p pd=0u as=82p ps=42u 
M1057 an3v0x2_0_a_24_8# an3v0x2_1_a an2v0x2_0_vss an2v0x2_0_vss nfet w=17u l=2u
+ ad=85p pd=44u as=0p ps=0u 
M1058 an3v0x2_0_a_31_8# an3v0x2_0_b an3v0x2_0_a_24_8# an2v0x2_0_vss nfet w=17u l=2u
+ ad=85p pd=44u as=0p ps=0u 
M1059 an3v0x2_0_zn an2v0x2_0_b an3v0x2_0_a_31_8# an2v0x2_0_vss nfet w=17u l=2u
+ ad=97p pd=48u as=0p ps=0u 
M1060 an3v0x2_2_vdd an2v0x2_0_zn nr3v0x2_0_a an3v0x2_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=166p ps=70u 
M1061 an2v0x2_0_zn an3v0x2_2_c an3v0x2_2_vdd an3v0x2_2_vdd pfet w=19u l=2u
+ ad=152p pd=54u as=0p ps=0u 
M1062 an3v0x2_2_vdd an2v0x2_0_b an2v0x2_0_zn an3v0x2_2_vdd pfet w=19u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1063 an2v0x2_0_vss an2v0x2_0_zn nr3v0x2_0_a an2v0x2_0_vss nfet w=14u l=2u
+ ad=0p pd=0u as=98p ps=42u 
M1064 an2v0x2_0_a_24_13# an3v0x2_2_c an2v0x2_0_vss an2v0x2_0_vss nfet w=13u l=2u
+ ad=65p pd=36u as=0p ps=0u 
M1065 an2v0x2_0_zn an2v0x2_0_b an2v0x2_0_a_24_13# an2v0x2_0_vss nfet w=13u l=2u
+ ad=77p pd=40u as=0p ps=0u 
M1066 nr2v0x2_0_a_11_39# an2v0x2_3_z an3v0x2_2_vdd an3v0x2_2_vdd pfet w=27u l=2u
+ ad=135p pd=64u as=0p ps=0u 
M1067 nd3v0x2_0_a an2v0x2_1_z nr2v0x2_0_a_11_39# an3v0x2_2_vdd pfet w=27u l=2u
+ ad=216p pd=70u as=0p ps=0u 
M1068 nr2v0x2_0_a_28_39# an2v0x2_1_z nd3v0x2_0_a an3v0x2_2_vdd pfet w=27u l=2u
+ ad=135p pd=64u as=0p ps=0u 
M1069 an3v0x2_2_vdd an2v0x2_3_z nr2v0x2_0_a_28_39# an3v0x2_2_vdd pfet w=27u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1070 nd3v0x2_0_a an2v0x2_3_z an2v0x2_0_vss an2v0x2_0_vss nfet w=15u l=2u
+ ad=120p pd=46u as=0p ps=0u 
M1071 an2v0x2_0_vss an2v0x2_1_z nd3v0x2_0_a an2v0x2_0_vss nfet w=15u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1072 an3v0x2_2_vdd or3v0x2_1_zn an2v0x2_3_b an3v0x2_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=166p ps=70u 
M1073 or3v0x2_1_a_24_38# an3v0x2_2_b an3v0x2_2_vdd an3v0x2_2_vdd pfet w=22u l=2u
+ ad=110p pd=54u as=0p ps=0u 
M1074 or3v0x2_1_a_31_38# an3v0x2_1_a or3v0x2_1_a_24_38# an3v0x2_2_vdd pfet w=22u l=2u
+ ad=110p pd=54u as=0p ps=0u 
M1075 or3v0x2_1_zn an3v0x2_2_a or3v0x2_1_a_31_38# an3v0x2_2_vdd pfet w=22u l=2u
+ ad=167p pd=60u as=0p ps=0u 
M1076 or3v0x2_1_a_48_38# an3v0x2_2_a or3v0x2_1_zn an3v0x2_2_vdd pfet w=19u l=2u
+ ad=95p pd=48u as=0p ps=0u 
M1077 or3v0x2_1_a_55_38# an3v0x2_1_a or3v0x2_1_a_48_38# an3v0x2_2_vdd pfet w=19u l=2u
+ ad=95p pd=48u as=0p ps=0u 
M1078 an3v0x2_2_vdd an3v0x2_2_b or3v0x2_1_a_55_38# an3v0x2_2_vdd pfet w=19u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1079 an2v0x2_0_vss or3v0x2_1_zn an2v0x2_3_b an2v0x2_0_vss nfet w=14u l=2u
+ ad=0p pd=0u as=98p ps=42u 
M1080 or3v0x2_1_zn an3v0x2_2_b an2v0x2_0_vss an2v0x2_0_vss nfet w=8u l=2u
+ ad=116p pd=62u as=0p ps=0u 
M1081 an2v0x2_0_vss an3v0x2_1_a or3v0x2_1_zn an2v0x2_0_vss nfet w=8u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1082 or3v0x2_1_zn an3v0x2_2_a an2v0x2_0_vss an2v0x2_0_vss nfet w=8u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1083 an3v0x2_2_vdd an2v0x2_1_zn an2v0x2_1_z an3v0x2_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=166p ps=70u 
M1084 an2v0x2_1_zn an2v0x2_4_z an3v0x2_2_vdd an3v0x2_2_vdd pfet w=19u l=2u
+ ad=152p pd=54u as=0p ps=0u 
M1085 an3v0x2_2_vdd an2v0x2_1_b an2v0x2_1_zn an3v0x2_2_vdd pfet w=19u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1086 an2v0x2_0_vss an2v0x2_1_zn an2v0x2_1_z an2v0x2_0_vss nfet w=14u l=2u
+ ad=0p pd=0u as=98p ps=42u 
M1087 an2v0x2_1_a_24_13# an2v0x2_4_z an2v0x2_0_vss an2v0x2_0_vss nfet w=13u l=2u
+ ad=65p pd=36u as=0p ps=0u 
M1088 an2v0x2_1_zn an2v0x2_1_b an2v0x2_1_a_24_13# an2v0x2_0_vss nfet w=13u l=2u
+ ad=77p pd=40u as=0p ps=0u 
M1089 an3v0x2_2_vdd an2v0x2_4_zn an2v0x2_4_z an3v0x2_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=166p ps=70u 
M1090 an2v0x2_4_zn an2v0x2_0_b an3v0x2_2_vdd an3v0x2_2_vdd pfet w=19u l=2u
+ ad=152p pd=54u as=0p ps=0u 
M1091 an3v0x2_2_vdd an3v0x2_2_b an2v0x2_4_zn an3v0x2_2_vdd pfet w=19u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1092 an2v0x2_0_vss an2v0x2_4_zn an2v0x2_4_z an2v0x2_0_vss nfet w=14u l=2u
+ ad=0p pd=0u as=98p ps=42u 
M1093 an2v0x2_4_a_24_13# an2v0x2_0_b an2v0x2_0_vss an2v0x2_0_vss nfet w=13u l=2u
+ ad=65p pd=36u as=0p ps=0u 
M1094 an2v0x2_4_zn an3v0x2_2_b an2v0x2_4_a_24_13# an2v0x2_0_vss nfet w=13u l=2u
+ ad=77p pd=40u as=0p ps=0u 
M1095 an3v0x2_2_b iv1v0x4_2_a an3v0x2_2_vdd an3v0x2_2_vdd pfet w=28u l=2u
+ ad=224p pd=72u as=0p ps=0u 
M1096 an3v0x2_2_vdd iv1v0x4_2_a an3v0x2_2_b an3v0x2_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1097 an3v0x2_2_b iv1v0x4_2_a an2v0x2_0_vss an2v0x2_0_vss nfet w=17u l=2u
+ ad=118p pd=50u as=0p ps=0u 
M1098 an2v0x2_0_vss iv1v0x4_2_a an3v0x2_2_b an2v0x2_0_vss nfet w=11u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1099 an3v0x2_2_vdd an2v0x2_3_zn an2v0x2_3_z an3v0x2_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=166p ps=70u 
M1100 an2v0x2_3_zn an2v0x2_2_z an3v0x2_2_vdd an3v0x2_2_vdd pfet w=19u l=2u
+ ad=152p pd=54u as=0p ps=0u 
M1101 an3v0x2_2_vdd an2v0x2_3_b an2v0x2_3_zn an3v0x2_2_vdd pfet w=19u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1102 an2v0x2_0_vss an2v0x2_3_zn an2v0x2_3_z an2v0x2_0_vss nfet w=14u l=2u
+ ad=0p pd=0u as=98p ps=42u 
M1103 an2v0x2_3_a_24_13# an2v0x2_2_z an2v0x2_0_vss an2v0x2_0_vss nfet w=13u l=2u
+ ad=65p pd=36u as=0p ps=0u 
M1104 an2v0x2_3_zn an2v0x2_3_b an2v0x2_3_a_24_13# an2v0x2_0_vss nfet w=13u l=2u
+ ad=77p pd=40u as=0p ps=0u 
M1105 an3v0x2_2_vdd an2v0x2_2_zn an2v0x2_2_z an3v0x2_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=166p ps=70u 
M1106 an2v0x2_2_zn an3v0x2_2_c an3v0x2_2_vdd an3v0x2_2_vdd pfet w=19u l=2u
+ ad=152p pd=54u as=0p ps=0u 
M1107 an3v0x2_2_vdd an3v0x2_0_b an2v0x2_2_zn an3v0x2_2_vdd pfet w=19u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1108 an2v0x2_0_vss an2v0x2_2_zn an2v0x2_2_z an2v0x2_0_vss nfet w=14u l=2u
+ ad=0p pd=0u as=98p ps=42u 
M1109 an2v0x2_2_a_24_13# an3v0x2_2_c an2v0x2_0_vss an2v0x2_0_vss nfet w=13u l=2u
+ ad=65p pd=36u as=0p ps=0u 
M1110 an2v0x2_2_zn an3v0x2_0_b an2v0x2_2_a_24_13# an2v0x2_0_vss nfet w=13u l=2u
+ ad=77p pd=40u as=0p ps=0u 
M1111 an3v0x2_2_vdd or3v0x2_0_zn an2v0x2_1_b an3v0x2_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=166p ps=70u 
M1112 or3v0x2_0_a_24_38# an3v0x2_0_b an3v0x2_2_vdd an3v0x2_2_vdd pfet w=22u l=2u
+ ad=110p pd=54u as=0p ps=0u 
M1113 or3v0x2_0_a_31_38# an3v0x2_2_a or3v0x2_0_a_24_38# an3v0x2_2_vdd pfet w=22u l=2u
+ ad=110p pd=54u as=0p ps=0u 
M1114 or3v0x2_0_zn an3v0x2_1_a or3v0x2_0_a_31_38# an3v0x2_2_vdd pfet w=22u l=2u
+ ad=167p pd=60u as=0p ps=0u 
M1115 or3v0x2_0_a_48_38# an3v0x2_1_a or3v0x2_0_zn an3v0x2_2_vdd pfet w=19u l=2u
+ ad=95p pd=48u as=0p ps=0u 
M1116 or3v0x2_0_a_55_38# an3v0x2_2_a or3v0x2_0_a_48_38# an3v0x2_2_vdd pfet w=19u l=2u
+ ad=95p pd=48u as=0p ps=0u 
M1117 an3v0x2_2_vdd an3v0x2_0_b or3v0x2_0_a_55_38# an3v0x2_2_vdd pfet w=19u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1118 an2v0x2_0_vss or3v0x2_0_zn an2v0x2_1_b an2v0x2_0_vss nfet w=14u l=2u
+ ad=0p pd=0u as=98p ps=42u 
M1119 or3v0x2_0_zn an3v0x2_0_b an2v0x2_0_vss an2v0x2_0_vss nfet w=8u l=2u
+ ad=116p pd=62u as=0p ps=0u 
M1120 an2v0x2_0_vss an3v0x2_2_a or3v0x2_0_zn an2v0x2_0_vss nfet w=8u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1121 or3v0x2_0_zn an3v0x2_1_a an2v0x2_0_vss an2v0x2_0_vss nfet w=8u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1122 an3v0x2_1_a iv1v0x4_1_a an3v0x2_2_vdd an3v0x2_2_vdd pfet w=28u l=2u
+ ad=224p pd=72u as=0p ps=0u 
M1123 an3v0x2_2_vdd iv1v0x4_1_a an3v0x2_1_a an3v0x2_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1124 an3v0x2_1_a iv1v0x4_1_a an2v0x2_0_vss an2v0x2_0_vss nfet w=17u l=2u
+ ad=118p pd=50u as=0p ps=0u 
M1125 an2v0x2_0_vss iv1v0x4_1_a an3v0x2_1_a an2v0x2_0_vss nfet w=11u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1126 an2v0x2_0_b iv1v0x4_0_a an3v0x2_2_vdd an3v0x2_2_vdd pfet w=28u l=2u
+ ad=224p pd=72u as=0p ps=0u 
M1127 an3v0x2_2_vdd iv1v0x4_0_a an2v0x2_0_b an3v0x2_2_vdd pfet w=28u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1128 an2v0x2_0_b iv1v0x4_0_a an2v0x2_0_vss an2v0x2_0_vss nfet w=17u l=2u
+ ad=118p pd=50u as=0p ps=0u 
M1129 an2v0x2_0_vss iv1v0x4_0_a an2v0x2_0_b an2v0x2_0_vss nfet w=11u l=2u
+ ad=0p pd=0u as=0p ps=0u 
C0 an2v0x2_1_z an2v0x2_0_vss 8.7fF
C1 an3v0x2_1_a or3v0x2_0_zn 4.1fF
C2 an2v0x2_0_vss or3v0x2_0_zn 10.9fF
C3 an3v0x2_2_zn an2v0x2_0_vss 8.8fF
C4 an2v0x2_3_zn an2v0x2_0_vss 8.9fF
C5 an3v0x2_2_vdd an3v0x2_1_zn 4.9fF
C6 an2v0x2_0_vss iv1v0x4_0_a 8.9fF
C7 an2v0x2_0_vss an3v0x2_2_z 10.7fF
C8 an3v0x2_2_a an3v0x2_2_vdd 41.3fF
C9 an3v0x2_2_vdd an2v0x2_4_zn 8.8fF
C10 an3v0x2_0_z an2v0x2_0_vss 36.9fF
C11 an3v0x2_2_zn an3v0x2_2_w_n4_32# 5.8fF
C12 an3v0x2_2_vdd an3v0x2_2_b 39.7fF
C13 an2v0x2_0_vss nr3v0x2_0_z 21.2fF
C14 an3v0x2_1_a an3v0x2_0_zn 2.5fF
C15 an2v0x2_0_vss an2v0x2_2_zn 8.9fF
C16 an3v0x2_1_a an2v0x2_0_b 2.5fF
C17 an2v0x2_0_vss an3v0x2_0_zn 8.8fF
C18 an2v0x2_0_vss an2v0x2_0_b 32.8fF
C19 an3v0x2_2_z an3v0x2_2_w_n4_32# 21.1fF
C20 an3v0x2_0_z an3v0x2_2_w_n4_32# 9.5fF
C21 an3v0x2_2_vdd iv1v0x4_1_a 9.9fF
C22 an2v0x2_0_vss nd3v0x2_0_c 18.9fF
C23 an3v0x2_2_vdd an2v0x2_2_z 9.4fF
C24 nr3v0x2_0_z an3v0x2_2_w_n4_32# 21.8fF
C25 an2v0x2_0_vss or3v0x2_1_zn 10.9fF
C26 an2v0x2_0_vss nd3v0x2_0_z 5.3fF
C27 an3v0x2_2_zn nr3v0x2_0_a 2.1fF
C28 an2v0x2_4_z an2v0x2_0_vss 9.8fF
C29 nd3v0x2_0_c an3v0x2_2_w_n4_32# 5.7fF
C30 an3v0x2_1_a an2v0x2_0_vss 57.3fF
C31 an3v0x2_0_b an2v0x2_0_vss 19.6fF
C32 an3v0x2_2_vdd an2v0x2_1_zn 8.8fF
C33 iv1v0x4_2_a an2v0x2_0_vss 8.9fF
C34 nd3v0x2_0_z an3v0x2_2_w_n4_32# 5.2fF
C35 an3v0x2_0_b an3v0x2_3_zn 3.6fF
C36 an2v0x2_1_z an3v0x2_2_vdd 22.0fF
C37 an2v0x2_0_vss an3v0x2_3_zn 8.8fF
C38 an3v0x2_1_a an3v0x2_2_w_n4_32# 8.3fF
C39 an2v0x2_0_vss nd3v0x2_0_a 21.1fF
C40 nr2v0x2_1_a nd3v0x2_0_c 3.8fF
C41 an2v0x2_0_vss an3v0x2_3_z 10.6fF
C42 an3v0x2_2_vdd or3v0x2_0_zn 9.0fF
C43 an2v0x2_0_vss an3v0x2_2_c 35.6fF
C44 an2v0x2_0_vss an2v0x2_1_b 5.9fF
C45 an3v0x2_2_vdd an3v0x2_2_zn 4.9fF
C46 an3v0x2_2_a or3v0x2_0_zn 3.3fF
C47 an3v0x2_2_vdd an2v0x2_3_zn 8.8fF
C48 nd3v0x2_0_a an3v0x2_2_w_n4_32# 6.2fF
C49 an3v0x2_2_vdd iv1v0x4_0_a 9.9fF
C50 an2v0x2_0_vss an2v0x2_0_zn 8.9fF
C51 an3v0x2_2_vdd an3v0x2_2_z 3.3fF
C52 an2v0x2_3_b an2v0x2_0_vss 15.0fF
C53 an3v0x2_0_z an3v0x2_2_vdd 2.3fF
C54 an2v0x2_0_vss nr2v0x2_1_a 22.9fF
C55 an3v0x2_2_c an3v0x2_2_w_n4_32# 11.6fF
C56 an3v0x2_2_vdd nr3v0x2_0_z 8.7fF
C57 an3v0x2_2_vdd an2v0x2_2_zn 8.8fF
C58 an2v0x2_0_vss nr3v0x2_0_a 19.9fF
C59 an2v0x2_3_z an2v0x2_0_vss 20.8fF
C60 an3v0x2_2_vdd an3v0x2_0_zn 10.7fF
C61 an3v0x2_2_vdd an2v0x2_0_b 49.9fF
C62 an3v0x2_2_a an3v0x2_0_zn 4.6fF
C63 an3v0x2_2_a an2v0x2_0_b 4.9fF
C64 an3v0x2_2_vdd nd3v0x2_0_c 5.0fF
C65 an3v0x2_2_b an2v0x2_0_b 2.5fF
C66 an3v0x2_2_vdd or3v0x2_1_zn 9.0fF
C67 nr3v0x2_0_a an3v0x2_2_w_n4_32# 15.0fF
C68 an3v0x2_2_vdd nd3v0x2_0_z 6.1fF
C69 an3v0x2_2_c nr3v0x2_0_a 2.5fF
C70 an2v0x2_4_z an3v0x2_2_vdd 10.7fF
C71 an3v0x2_1_a an3v0x2_2_vdd 72.4fF
C72 an3v0x2_1_zn an2v0x2_0_vss 8.8fF
C73 an3v0x2_0_b an3v0x2_2_vdd 47.7fF
C74 an3v0x2_2_a an3v0x2_1_a 6.8fF
C75 iv1v0x4_2_a an3v0x2_2_vdd 9.9fF
C76 an3v0x2_2_a an2v0x2_0_vss 61.9fF
C77 an3v0x2_1_a an3v0x2_2_b 5.2fF
C78 an2v0x2_4_zn an2v0x2_0_vss 8.9fF
C79 an3v0x2_2_a iv1v0x4_2_a 2.2fF
C80 an3v0x2_2_b an2v0x2_0_vss 23.0fF
C81 an3v0x2_2_vdd an3v0x2_3_zn 10.7fF
C82 an3v0x2_1_zn an3v0x2_2_w_n4_32# 5.8fF
C83 an3v0x2_2_vdd nd3v0x2_0_a 9.6fF
C84 an3v0x2_2_vdd an3v0x2_2_w_n4_32# 87.6fF
C85 an3v0x2_2_vdd an3v0x2_3_z 15.4fF
C86 an3v0x2_2_a an3v0x2_2_w_n4_32# 8.1fF
C87 an2v0x2_0_vss iv1v0x4_1_a 8.9fF
C88 an3v0x2_2_vdd an2v0x2_1_b 14.2fF
C89 an3v0x2_2_vdd an3v0x2_2_c 23.8fF
C90 an2v0x2_0_vss an2v0x2_2_z 11.1fF
C91 an3v0x2_2_b an3v0x2_2_w_n4_32# 21.4fF
C92 an3v0x2_2_a an2v0x2_1_b 2.2fF
C93 an3v0x2_2_vdd an2v0x2_0_zn 8.8fF
C94 an3v0x2_2_vdd an2v0x2_3_b 13.7fF
C95 an3v0x2_2_vdd nr2v0x2_1_a 7.1fF
C96 an2v0x2_1_zn an2v0x2_0_vss 8.9fF
C97 an3v0x2_2_vdd nr3v0x2_0_a 4.0fF
C98 an2v0x2_3_z an3v0x2_2_vdd 9.1fF
C99 an3v0x2_2_c 0 18.7fF
C100 an3v0x2_2_vdd 0 379.0fF
C101 an2v0x2_0_vss 0 10.8fF
C102 nr3v0x2_0_a 0 8.6fF

v_dd an3v0x2_2_vdd 0 5
v_ss an2v0x2_0_vss 0 0
v_gg_f iv1v0x4_1_a 0 PULSE(5 0 0 0.1n 0.1n 150n 300n)
v_gg_e iv1v0x4_2_a 0 PULSE(5 0 0 0.1n 0.1n 300n 600n)
v_gg_d iv1v0x4_0_a 0 PULSE(5 0 0 0.1n 0.1n 600n 1200n)
v_gg_c an3v0x2_2_a 0 PULSE(5 0 0 0.1n 0.1n 1200n 2400n)
v_gg_b an3v0x2_0_b 0 PULSE(5 0 0 0.1n 0.1n 2400n 4800n)
v_gg_a an3v0x2_2_c 0 PULSE(5 0 0 0.1n 0.1n 4800n 9600n)

.control
 tran 1n 9600n
 plot (an3v0x2_2_c + 5) (an3v0x2_0_b) (an3v0x2_2_a - 5) (iv1v0x4_0_a - 10) (iv1v0x4_2_a - 15) (iv1v0x4_1_a - 20) ( nd3v0x2_0_z - 25)
.endc

.end