* Spice description of oai22_x2
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:10
*
.subckt oai22_x2 a1 a2 b1 b2 vdd vss z 
M1b n1b   a1    vdd   vdd p  L=0.13U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U   
M2b z     a2    n1b   vdd p  L=0.13U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U   
M2a sig6  a2    z     vdd p  L=0.13U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U   
M1a vdd   a1    sig6  vdd p  L=0.13U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U   
M3b n2b   b1    vdd   vdd p  L=0.13U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U   
M4a n2a   b2    z     vdd p  L=0.13U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U   
M3a vdd   b1    n2a   vdd p  L=0.13U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U   
M4b z     b2    n2b   vdd p  L=0.13U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U   
M8  z     b2    sig1  vss n  L=0.13U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U  
M7  sig1  b1    z     vss n  L=0.13U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U  
M6  sig1  a2    vss   vss n  L=0.13U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U  
M5  vss   a1    sig1  vss n  L=0.13U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U  
C12 a2    vss   1.379f
C10 b1    vss   2.045f
C9  a1    vss   2.268f
C8  b2    vss   1.050f
C5  vdd   vss   2.618f
C2  z     vss   4.620f
C1  sig1  vss   0.918f
.ends
