* Tue Aug 10 11:21:07 CEST 2004
.subckt oai22_x1 a1 a2 b1 b2 vdd vss z 
*SPICE circuit <oai22_x1> from XCircuit v3.10

m1 z b1 n2 vss n w=17u l=2.3636u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m2 int14 b1 vdd vdd p w=39u l=2.3636u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m3 n1 a1 vdd vdd p w=39u l=2.3636u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m4 z b2 int14 vdd p w=39u l=2.3636u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m5 n2 a2 vss vss n w=17u l=2.3636u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m6 n2 a1 vss vss n w=17u l=2.3636u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m7 z b2 n2 vss n w=17u l=2.3636u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m8 z a2 n1 vdd p w=39u l=2.3636u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
.ends
