* Thu Jan 11 12:49:18 CET 2007
.subckt iv1v0x12 a vdd vss z
*SPICE circuit <iv1v0x12> from XCircuit v3.20

m1 z a vss vss n w=120u l=2u ad='120u*5u+12p' as='120u*5u+12p' pd='120u*2+14u' ps='120u*2+14u'
m2 z a vdd vdd p w=168u l=2u ad='168u*5u+12p' as='168u*5u+12p' pd='168u*2+14u' ps='168u*2+14u'
.ends
