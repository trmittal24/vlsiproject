* Spice description of vfeed8
* Spice driver version 134999461
* Date 17/05/2007 at  9:36:29
* wsclib 0.13um values
.subckt vfeed8 vdd vss
.ends
