* Tue Apr  4 18:58:27 CEST 2006
.subckt iv1v3x1 a vdd vss z 
*SPICE circuit <iv1v3x1> from XCircuit v3.20

m1 z a vss vss n w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m2 z a vdd vdd p w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
.ends
