magic
tech scmos
timestamp 1523087730
<< metal1 >>
rect -15 71 -12 75
rect -4 68 6 76
rect 29 68 36 76
rect 94 68 100 76
rect -15 50 -12 54
rect 177 44 180 48
rect -15 26 -12 30
rect -6 4 4 12
rect 29 4 36 12
rect 94 4 100 12
<< metal2 >>
rect -13 71 -12 74
rect -8 71 83 74
rect -8 50 24 54
rect 79 47 83 71
rect 148 54 171 58
rect 148 48 152 54
rect 107 44 152 48
rect 6 30 10 36
rect 157 39 161 46
rect 167 48 171 54
rect 167 44 173 48
rect 42 36 161 39
rect 38 35 161 36
rect 6 26 79 30
rect -12 22 -8 26
rect 150 22 154 26
rect -12 18 154 22
<< m2contact >>
rect -12 71 -8 75
rect -12 50 -8 54
rect 24 50 28 54
rect 79 43 83 47
rect 103 44 107 48
rect 157 46 161 50
rect 173 44 177 48
rect 6 36 10 40
rect 38 36 42 40
rect -12 26 -8 30
rect 79 26 83 30
rect 150 26 154 30
use /home/dipanshu/Desktop/vlsiproject/pharosc_8.4/magic/cells/vsclib/iv1v0x2  iv1v0x2_0
timestamp 1523087564
transform 1 0 4 0 1 4
box -4 -4 28 76
use /home/dipanshu/Desktop/vlsiproject/pharosc_8.4/magic/cells/vsclib/an2v0x3  an2v0x3_0
timestamp 1523087564
transform 1 0 36 0 1 4
box -4 -4 60 76
use /home/dipanshu/Desktop/vlsiproject/pharosc_8.4/magic/cells/vsclib/or2v0x3  or2v0x3_0
timestamp 1523087564
transform 1 0 100 0 1 4
box -4 -4 68 76
<< labels >>
rlabel metal1 -13 52 -13 52 3 b
rlabel metal1 -14 73 -14 73 3 c
rlabel metal1 -13 28 -13 28 3 a
rlabel metal1 -4 8 -4 8 1 gnd
rlabel metal1 -3 69 -3 69 1 vdd
rlabel metal1 178 45 178 45 7 out
<< end >>
