* Mon Aug 16 14:11:00 CEST 2004
.subckt nr4v0x1 a b c d vdd vss z 
*SPICE circuit <nr4v0x1> from XCircuit v3.10

m1 z a vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m2 z b vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m3 z d vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m4 n1 a vdd vdd p w=43u l=2u ad='43u*5u+12p' as='43u*5u+12p' pd='43u*2+14u' ps='43u*2+14u'
m5 n2 b n1 vdd p w=43u l=2u ad='43u*5u+12p' as='43u*5u+12p' pd='43u*2+14u' ps='43u*2+14u'
m6 n3 c n2 vdd p w=43u l=2u ad='43u*5u+12p' as='43u*5u+12p' pd='43u*2+14u' ps='43u*2+14u'
m7 z c vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m8 z d n3 vdd p w=43u l=2u ad='43u*5u+12p' as='43u*5u+12p' pd='43u*2+14u' ps='43u*2+14u'
.ends
