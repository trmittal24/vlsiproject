* Spice description of aoi22_x05
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:09
*
.subckt aoi22_x05 a1 a2 b1 b2 vdd vss z 
M2  vdd   a2    2     vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M1  2     a1    z     vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M3  z     b1    2     vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M4  2     b2    vdd   vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M5  n2    a1    vss   vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M6  vss   a2    sig1  vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M8  sig1  b2    z     vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M7  z     b1    n2    vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
C10 2     vss   0.918f
C9  vdd   vss   1.290f
C8  b1    vss   1.383f
C7  b2    vss   1.623f
C6  a1    vss   1.409f
C5  a2    vss   1.661f
C4  z     vss   2.505f
.ends
