* Spice description of oai22_x05
* Spice driver version 134999461
* Date 31/05/2007 at 21:35:18
* vxlib 0.13um values
.subckt oai22_x05 a1 a2 b1 b2 vdd vss z
M1  n1    a1    vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M2  z     a2    n1    vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M3  vdd   b1    3     vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M4  3     b2    z     vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M5  n3    a1    vss   vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M6  vss   a2    n3    vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M7  z     b1    n3    vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M8  n3    b2    z     vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
C6  a1    vss   0.594f
C5  a2    vss   0.757f
C7  b1    vss   0.591f
C4  b2    vss   0.614f
C2  n3    vss   0.526f
C3  z     vss   0.927f
.ends
