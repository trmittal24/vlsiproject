* Spice description of nd2av0x1
* Spice driver version 134999461
* Date 17/05/2007 at  9:17:13
* wsclib 0.13um values
.subckt nd2av0x1 a b vdd vss z
M01 06    a     vdd   vdd p  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
M02 06    a     vss   vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M03 z     b     vdd   vdd p  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
M04 sig3  b     z     vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M05 vdd   06    z     vdd p  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
M06 vss   06    sig3  vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
C5  06    vss   0.570f
C6  a     vss   0.465f
C4  b     vss   0.515f
C2  z     vss   0.590f
.ends
