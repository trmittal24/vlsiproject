* Spice description of an3_x2
* Spice driver version 134999461
* Date 31/05/2007 at 21:32:21
* vxlib 0.13um values
.subckt an3_x2 a b c vdd vss z
M1a zn    a     vdd   vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M1b vdd   b     zn    vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M1c zn    c     vdd   vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M1z vdd   zn    z     vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M2a vss   a     sig5  vss n  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M2b sig5  b     sig4  vss n  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M2c sig4  c     zn    vss n  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M2z z     zn    vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
C9  a     vss   0.649f
C8  b     vss   0.649f
C7  c     vss   0.677f
C1  z     vss   0.891f
C3  zn    vss   1.125f
.ends
