* Sat Aug 27 22:10:09 CEST 2005
.subckt iv1v4x8 a vdd vss z 
*SPICE circuit <iv1v4x8> from XCircuit v3.20

m1 z a vss vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m2 z a vdd vdd p w=128u l=2u ad='128u*5u+12p' as='128u*5u+12p' pd='128u*2+14u' ps='128u*2+14u'
.ends
