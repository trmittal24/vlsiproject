* Tue Aug 10 11:21:07 CEST 2004
.subckt iv1_x8 a vdd vss z 
*SPICE circuit <iv1_x8> from XCircuit v3.10

m1 z a vss vss n w=72u l=2u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
m2 z a vdd vdd p w=145u l=2u ad='145u*5u+12p' as='145u*5u+12p' pd='145u*2+14u' ps='145u*2+14u'
.ends
