* Sat Apr  9 11:31:04 CEST 2005
.subckt nr3v0x3 a b c vdd vss z 
*SPICE circuit <nr3v0x3> from XCircuit v3.20

m1 z a vss vss n w=19u l=2u ad='19u*5u+12p' as='19u*5u+12p' pd='19u*2+14u' ps='19u*2+14u'
m2 z c vss vss n w=19u l=2u ad='19u*5u+12p' as='19u*5u+12p' pd='19u*2+14u' ps='19u*2+14u'
m3 n1 a vdd vdd p w=104u l=2u ad='104u*5u+12p' as='104u*5u+12p' pd='104u*2+14u' ps='104u*2+14u'
m4 n2 b n1 vdd p w=104u l=2u ad='104u*5u+12p' as='104u*5u+12p' pd='104u*2+14u' ps='104u*2+14u'
m5 z b vss vss n w=19u l=2u ad='19u*5u+12p' as='19u*5u+12p' pd='19u*2+14u' ps='19u*2+14u'
m6 z c n2 vdd p w=104u l=2u ad='104u*5u+12p' as='104u*5u+12p' pd='104u*2+14u' ps='104u*2+14u'
.ends
