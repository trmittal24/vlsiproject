* Spice description of o2_x4
* Spice driver version 134999461
* Date 21/07/2007 at 19:31:31
* sxlib 0.13um values
.subckt o2_x4 i0 i1 q vdd vss
Mtr_00001 q     sig1  vss   vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00002 sig1  i0    vss   vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00003 vss   i1    sig1  vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00004 vss   sig1  q     vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00005 sig5  i1    sig1  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00006 vdd   i0    sig5  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00007 q     sig1  vdd   vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00008 vdd   sig1  q     vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
C6  i0    vss   0.908f
C7  i1    vss   0.668f
C3  q     vss   0.883f
C1  sig1  vss   0.865f
.ends
