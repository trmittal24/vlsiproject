* Wed Apr 11 09:12:53 CEST 2007
.subckt xor2v0x4 a b vdd vss z
*SPICE circuit <xor2v0x4> from XCircuit v3.4 rev 26

m1 z bn an vdd p w=75u l=2u ad='75u*5u+12p' as='75u*5u+12p' pd='75u*2+14u' ps='75u*2+14u'
m2 bn b vss vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m3 an a vss vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m4 z an n1 vss n w=48u l=2u ad='48u*5u+12p' as='48u*5u+12p' pd='48u*2+14u' ps='48u*2+14u'
m5 n1 bn vss vss n w=48u l=2u ad='48u*5u+12p' as='48u*5u+12p' pd='48u*2+14u' ps='48u*2+14u'
m6 an a vdd vdd p w=75u l=2u ad='75u*5u+12p' as='75u*5u+12p' pd='75u*2+14u' ps='75u*2+14u'
m7 bn b vdd vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
m8 z b an vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m9 z an bn vdd p w=113u l=2u ad='113u*5u+12p' as='113u*5u+12p' pd='113u*2+14u' ps='113u*2+14u'
.ends
