* Spice description of iv1_x2
* Spice driver version 134999461
* Date 31/05/2007 at 21:33:54
* vxlib 0.13um values
.subckt iv1_x2 a vdd vss z
M1  vdd   a     z     vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M2  z     a     vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
C4  a     vss   0.439f
C2  z     vss   0.778f
.ends
