* Sat Apr  9 10:46:06 CEST 2005
.subckt nd2av0x8 a b vdd vss z 
*SPICE circuit <nd2av0x8> from XCircuit v3.20

m1 an a vss vss n w=22u l=2u ad='22u*5u+12p' as='22u*5u+12p' pd='22u*2+14u' ps='22u*2+14u'
m2 n1 b vss vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m3 an a vdd vdd p w=44u l=2u ad='44u*5u+12p' as='44u*5u+12p' pd='44u*2+14u' ps='44u*2+14u'
m4 z b vdd vdd p w=96u l=2u ad='96u*5u+12p' as='96u*5u+12p' pd='96u*2+14u' ps='96u*2+14u'
m5 z an n1 vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m6 z an vdd vdd p w=96u l=2u ad='96u*5u+12p' as='96u*5u+12p' pd='96u*2+14u' ps='96u*2+14u'
.ends
