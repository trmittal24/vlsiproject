* Sat Aug 27 19:34:35 CEST 2005
.subckt nd2v4x6 a b vdd vss z 
*SPICE circuit <nd2v4x6> from XCircuit v3.20

m1 n1 a vss vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m2 z a vdd vdd p w=91u l=2u ad='91u*5u+12p' as='91u*5u+12p' pd='91u*2+14u' ps='91u*2+14u'
m3 z b n1 vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m4 z b vdd vdd p w=91u l=2u ad='91u*5u+12p' as='91u*5u+12p' pd='91u*2+14u' ps='91u*2+14u'
.ends
