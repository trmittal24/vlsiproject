* Sun Nov 28 16:58:20 CET 2004
.subckt nd2abv0x05 a b vdd vss z 
*SPICE circuit <nd2abv0x05> from XCircuit v3.20

m1 bn b vss vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m2 an a vss vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m3 bn b vdd vdd p w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m4 an a vdd vdd p w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m5 n1 an vss vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m6 z an vdd vdd p w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m7 z bn n1 vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m8 z bn vdd vdd p w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
.ends
