* Spice description of nd2a_x2
* Spice driver version 134999461
* Date 31/05/2007 at 21:34:18
* vxlib 0.13um values
.subckt nd2a_x2 a b vdd vss z
M1a sig3  a     vdd   vdd p  L=0.12U  W=1.65U  AS=0.43725P  AD=0.43725P  PS=3.83U   PD=3.83U
M1  z     b     vdd   vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M2a vss   a     sig3  vss n  L=0.12U  W=0.825U AS=0.218625P AD=0.218625P PS=2.18U   PD=2.18U
M2  vdd   sig3  z     vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M3  z     b     sig1  vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M4  sig1  sig3  vss   vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
C7  a     vss   0.640f
C6  b     vss   0.574f
C3  sig3  vss   0.727f
C4  z     vss   0.891f
.ends
