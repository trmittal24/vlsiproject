* Spice description of bf1_y05
* Spice driver version 134999461
* Date 22/07/2007 at 10:57:50
* vsxlib 0.13um values
.subckt bf1_y05 a vdd vss z
M1a 2z    a     vdd   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M1z vdd   2z    z     vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M2a vss   a     2z    vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M2z z     2z    vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
C4  2z    vss   0.699f
C3  a     vss   0.490f
C2  z     vss   0.520f
.ends
