* Wed Apr 11 09:50:31 CEST 2007
.subckt xor2v0x6 a b vdd vss z
*SPICE circuit <xor2v0x6> from XCircuit v3.4 rev 26

m1 z bn an vdd p w=109u l=2u ad='109u*5u+12p' as='109u*5u+12p' pd='109u*2+14u' ps='109u*2+14u'
m2 bn b vss vss n w=54u l=2u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m3 an a vss vss n w=54u l=2u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m4 z an n1 vss n w=72u l=2u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
m5 n1 bn vss vss n w=72u l=2u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
m6 an a vdd vdd p w=108u l=2u ad='108u*5u+12p' as='108u*5u+12p' pd='108u*2+14u' ps='108u*2+14u'
m7 bn b vdd vdd p w=162u l=2u ad='162u*5u+12p' as='162u*5u+12p' pd='162u*2+14u' ps='162u*2+14u'
m8 z b an vss n w=54u l=2u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m9 z an bn vdd p w=162u l=2u ad='162u*5u+12p' as='162u*5u+12p' pd='162u*2+14u' ps='162u*2+14u'
.ends
