* Tue Aug 10 11:21:07 CEST 2004
.subckt iv1_y2 a vdd vss z 
*SPICE circuit <iv1_y2> from XCircuit v3.10

m1 z a vss vss n w=16u l=2u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m2 z a vdd vdd p w=36u l=2u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
.ends
