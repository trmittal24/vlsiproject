* Spice description of aon21bv0x05
* Spice driver version 134999461
* Date 17/05/2007 at  9:03:09
* vsclib 0.13um values
.subckt aon21bv0x05 a1 a2 b vdd vss z
M01 vdd   a2    08    vdd p  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M02 08    a2    n1    vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M03 08    a1    vdd   vdd p  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M04 n1    a1    vss   vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M05 z     b     vdd   vdd p  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M06 n2    b     z     vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M07 vdd   08    z     vdd p  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M08 vss   08    n2    vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
C6  08    vss   0.583f
C4  a1    vss   0.433f
C8  a2    vss   0.582f
C5  b     vss   0.461f
C1  z     vss   0.634f
.ends
