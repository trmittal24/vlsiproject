* Spice description of vfeed8
* Spice driver version 134999461
* Date 22/07/2007 at 11:00:30
* vsxlib 0.13um values
.subckt vfeed8 vdd vss
.ends
