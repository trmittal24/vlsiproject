* Spice description of nr2a_x1
* Spice driver version 134999461
* Date 22/07/2007 at 10:59:23
* vsxlib 0.13um values
.subckt nr2a_x1 a b vdd vss z
M1a 3z    a     vdd   vdd p  L=0.12U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U
M1z vdd   3z    2z    vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M2a vss   a     3z    vss n  L=0.12U  W=0.605U AS=0.160325P AD=0.160325P PS=1.74U   PD=1.74U
M2z 2z    b     z     vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M3z z     3z    vss   vss n  L=0.12U  W=0.605U AS=0.160325P AD=0.160325P PS=1.74U   PD=1.74U
M4z vss   b     z     vss n  L=0.12U  W=0.605U AS=0.160325P AD=0.160325P PS=1.74U   PD=1.74U
C4  3z    vss   0.619f
C5  a     vss   0.653f
C3  b     vss   0.692f
C1  z     vss   0.763f
.ends
