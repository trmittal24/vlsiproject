* Tue Aug 10 11:21:08 CEST 2004
.subckt xnr2_x1 a b vdd vss z 
*SPICE circuit <xnr2_x1> from XCircuit v3.10

m1 bn b vdd vdd p w=37u l=2u ad='37u*5u+12p' as='37u*5u+12p' pd='37u*2+14u' ps='37u*2+14u'
m2 z bn n1 vdd p w=37u l=2u ad='37u*5u+12p' as='37u*5u+12p' pd='37u*2+14u' ps='37u*2+14u'
m3 z b an vdd p w=37u l=2u ad='37u*5u+12p' as='37u*5u+12p' pd='37u*2+14u' ps='37u*2+14u'
m4 bn b vss vss n w=16u l=2u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m5 an a vss vss n w=16u l=2u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m6 z an bn vss n w=16u l=2u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m7 an a vdd vdd p w=37u l=2u ad='37u*5u+12p' as='37u*5u+12p' pd='37u*2+14u' ps='37u*2+14u'
m8 z bn an vss n w=16u l=2u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m9 n1 an vdd vdd p w=37u l=2u ad='37u*5u+12p' as='37u*5u+12p' pd='37u*2+14u' ps='37u*2+14u'
.ends
