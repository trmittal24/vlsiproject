* Spice description of powmid_x0
* Spice driver version 134999461
* Date 22/07/2007 at 11:00:09
* vsxlib 0.13um values
.subckt powmid_x0 vdd vss
.ends
