* Spice description of aoi21_x1
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:09
*
.subckt aoi21_x1 a1 a2 b vdd vss z 
M2  n2    a2    vdd   vdd p  L=0.13U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U  
M3  z     b     n2    vdd p  L=0.13U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U  
M1  vdd   a1    n2    vdd p  L=0.13U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U  
M6  z     b     vss   vss n  L=0.13U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U  
M5  sig3  a2    z     vss n  L=0.13U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U   
M4  vss   a1    sig3  vss n  L=0.13U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U   
C8  a2    vss   0.979f
C7  a1    vss   0.964f
C6  b     vss   1.613f
C5  vdd   vss   1.003f
C4  n2    vss   0.529f
C1  z     vss   2.253f
.ends
