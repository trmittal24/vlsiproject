* Mon Aug 16 14:22:57 CEST 2004
.subckt noa22_x1 i0 i1 i2 nq vdd vss 
*SPICE circuit <noa22_x1> from XCircuit v3.10

m1 nq i1 n1 vdd p w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m2 n1 i2 vdd vdd p w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m3 n2 i0 vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m4 nq i2 vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m5 nq i1 n2 vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m6 nq i0 n1 vdd p w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
.ends
