* Tue Aug 10 21:18:16 CEST 2004
.subckt ha2_x2 a b co so vdd vss 
*SPICE circuit <ha2_x2> from XCircuit v3.10

m1 so son vss vss n w=19u l=2u ad='19u*5u+12p' as='19u*5u+12p' pd='19u*2+14u' ps='19u*2+14u'
m2 son a n2 vss n w=15u l=2u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m3 so son vdd vdd p w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m4 son vss vdd vdd p w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m5 co vss vss vss n w=19u l=2u ad='19u*5u+12p' as='19u*5u+12p' pd='19u*2+14u' ps='19u*2+14u'
m6 co vss vdd vdd p w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m7 n3 a vdd vdd p w=34u l=2u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
m8 son b n3 vdd p w=34u l=2u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
m9 n2 vss vss vss n w=15u l=2u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m10 son b n2 vss n w=15u l=2u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m11 n1 b vss vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m12 vss b vdd vdd p w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m13 vss a vdd vdd p w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m14 vss a n1 vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
.ends
