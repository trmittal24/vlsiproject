* Spice description of nd2_x05
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:10
*
.subckt nd2_x05 a b vdd vss z 
M1  z     b     vdd   vdd p  L=0.13U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U  
M2  vdd   a     z     vdd p  L=0.13U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U  
M4  sig3  a     vss   vss n  L=0.13U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U  
M3  z     b     sig3  vss n  L=0.13U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U  
C6  a     vss   1.023f
C5  b     vss   1.075f
C4  vdd   vss   1.273f
C2  z     vss   1.712f
.ends
