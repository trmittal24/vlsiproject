* Spice description of nr2_x05
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:10
*
.subckt nr2_x05 a b vdd vss z 
M2  vdd   a     sig3  vdd p  L=0.13U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U  
M1  sig3  b     z     vdd p  L=0.13U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U  
M3  vss   b     z     vss n  L=0.13U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U  
M4  z     a     vss   vss n  L=0.13U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U  
C6  a     vss   0.979f
C5  b     vss   0.991f
C4  vdd   vss   1.078f
C1  z     vss   1.920f
.ends
