* Tue Aug 10 11:21:07 CEST 2004
.subckt nd2_x2 a b vdd vss z 
*SPICE circuit <nd2_x2> from XCircuit v3.10

m1 n1 a vss vss n w=33u l=2u ad='33u*5u+12p' as='33u*5u+12p' pd='33u*2+14u' ps='33u*2+14u'
m2 z a vdd vdd p w=39u l=2u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m3 z b n1 vss n w=33u l=2u ad='33u*5u+12p' as='33u*5u+12p' pd='33u*2+14u' ps='33u*2+14u'
m4 z b vdd vdd p w=39u l=2u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
.ends
