* Sun Dec 18 19:34:49 CET 2005
.subckt iv1v1x8 a vdd vss z 
*SPICE circuit <iv1v1x8> from XCircuit v3.20

m1 z a vss vss n w=69u l=2u ad='69u*5u+12p' as='69u*5u+12p' pd='69u*2+14u' ps='69u*2+14u'
m2 z a vdd vdd p w=104u l=2u ad='104u*5u+12p' as='104u*5u+12p' pd='104u*2+14u' ps='104u*2+14u'
.ends
