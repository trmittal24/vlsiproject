* Spice description of nd2_x2
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:10
*
.subckt nd2_x2 a b vdd vss z 
M1  z     b     vdd   vdd p  L=0.13U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U  
M2  vdd   a     z     vdd p  L=0.13U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U  
M3  z     b     sig1  vss n  L=0.13U  W=1.76U  AS=0.4664P   AD=0.4664P   PS=4.05U   PD=4.05U  
M4  sig1  a     vss   vss n  L=0.13U  W=1.76U  AS=0.4664P   AD=0.4664P   PS=4.05U   PD=4.05U  
C6  a     vss   0.926f
C5  b     vss   0.966f
C4  vdd   vss   1.273f
C3  z     vss   2.487f
.ends
