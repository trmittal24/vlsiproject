* Sun Apr  9 08:49:38 CEST 2006
.subckt oai21v0x6 a1 a2 b vdd vss z 
*SPICE circuit <oai21v0x6> from XCircuit v3.20

m1 n2 a1 vdd vdd p w=160u l=2.3636u ad='160u*5u+12p' as='160u*5u+12p' pd='160u*2+14u' ps='160u*2+14u'
m2 z b vdd vdd p w=84u l=2.3636u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m3 n1 a2 vss vss n w=70u l=2.3636u ad='70u*5u+12p' as='70u*5u+12p' pd='70u*2+14u' ps='70u*2+14u'
m4 n1 a1 vss vss n w=70u l=2.3636u ad='70u*5u+12p' as='70u*5u+12p' pd='70u*2+14u' ps='70u*2+14u'
m5 z b n1 vss n w=70u l=2.3636u ad='70u*5u+12p' as='70u*5u+12p' pd='70u*2+14u' ps='70u*2+14u'
m6 z a2 n2 vdd p w=160u l=2.3636u ad='160u*5u+12p' as='160u*5u+12p' pd='160u*2+14u' ps='160u*2+14u'
.ends
