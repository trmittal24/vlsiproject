* Mon Aug 16 14:11:01 CEST 2004
.subckt oai22v0x2 a1 a2 b1 b2 vdd vss z 
*SPICE circuit <oai22v0x2> from XCircuit v3.10

m1 z b1 n2 vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m2 int14 b1 vdd vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m3 n1 a1 vdd vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m4 z b2 int14 vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m5 n2 a2 vss vss n w=23u l=2u ad='23u*5u+12p' as='23u*5u+12p' pd='23u*2+14u' ps='23u*2+14u'
m6 n2 a1 vss vss n w=23u l=2u ad='23u*5u+12p' as='23u*5u+12p' pd='23u*2+14u' ps='23u*2+14u'
m7 z b2 n2 vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m8 z a2 n1 vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
.ends
