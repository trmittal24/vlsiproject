* Mon Aug 16 14:10:58 CEST 2004
.subckt nd2abv0x3 a b vdd vss z 
*SPICE circuit <nd2abv0x3> from XCircuit v3.10

m1 bn b vss vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m2 an a vss vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m3 bn b vdd vdd p w=26u l=2.3636u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m4 an a vdd vdd p w=26u l=2.3636u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m5 n1 an vss vss n w=36u l=2.3636u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
m6 z an vdd vdd p w=44u l=2.3636u ad='44u*5u+12p' as='44u*5u+12p' pd='44u*2+14u' ps='44u*2+14u'
m7 z bn n1 vss n w=36u l=2.3636u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
m8 z bn vdd vdd p w=44u l=2.3636u ad='44u*5u+12p' as='44u*5u+12p' pd='44u*2+14u' ps='44u*2+14u'
.ends
