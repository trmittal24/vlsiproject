* Sun Apr  2 21:56:03 CEST 2006
.subckt nd2v3x3 a b vdd vss z 
*SPICE circuit <nd2v3x3> from XCircuit v3.20

m1 n1 a vss vss n w=57u l=2u ad='57u*5u+12p' as='57u*5u+12p' pd='57u*2+14u' ps='57u*2+14u'
m2 z a vdd vdd p w=34u l=2u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
m3 z b n1 vss n w=57u l=2u ad='57u*5u+12p' as='57u*5u+12p' pd='57u*2+14u' ps='57u*2+14u'
m4 z b vdd vdd p w=34u l=2u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
.ends
