* Sun Apr  9 08:49:34 CEST 2006
.subckt oai21v0x3 a1 a2 b vdd vss z 
*SPICE circuit <oai21v0x3> from XCircuit v3.20

m1 n2 a1 vdd vdd p w=75u l=2.3636u ad='75u*5u+12p' as='75u*5u+12p' pd='75u*2+14u' ps='75u*2+14u'
m2 z b vdd vdd p w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m3 n1 a2 vss vss n w=34u l=2.3636u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
m4 n1 a1 vss vss n w=34u l=2.3636u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
m5 z b n1 vss n w=34u l=2.3636u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
m6 z a2 n2 vdd p w=75u l=2.3636u ad='75u*5u+12p' as='75u*5u+12p' pd='75u*2+14u' ps='75u*2+14u'
.ends
