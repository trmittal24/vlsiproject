* Spice description of nd2v0x2
* Spice driver version 134999461
* Date  6/02/2007 at 12:03:11
* rgalib 0.13um values
.subckt nd2v0x2 a b vdd vss z
Mtr_00001 sig3  a     vss   vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00002 z     b     sig3  vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00003 z     a     vdd   vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
Mtr_00004 vdd   b     z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
C4  a     vss   0.408f
C5  b     vss   0.408f
C2  z     vss   0.707f
.ends
