* Spice description of bf1_x2
* Spice driver version 134999461
* Date 31/05/2007 at 21:33:03
* vxlib 0.13um values
.subckt bf1_x2 a vdd vss z
M1a an    a     vdd   vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
M1z vdd   an    z     vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M2a vss   a     an    vss n  L=0.12U  W=0.715U AS=0.189475P AD=0.189475P PS=1.96U   PD=1.96U
M2z z     an    vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
C5  a     vss   0.457f
C3  an    vss   0.751f
C1  z     vss   0.677f
.ends
