* Mon Aug 16 14:10:58 CEST 2004
.subckt iv1v0x6 a vdd vss z 
*SPICE circuit <iv1v0x6> from XCircuit v3.10

m1 z a vss vss n w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m2 z a vdd vdd p w=81u l=2u ad='81u*5u+12p' as='81u*5u+12p' pd='81u*2+14u' ps='81u*2+14u'
.ends
