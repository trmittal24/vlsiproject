* Sat Aug 27 22:10:27 CEST 2005
.subckt iv1v5x1 a vdd vss z 
*SPICE circuit <iv1v5x1> from XCircuit v3.20

m1 z a vss vss n w=7u l=2.3636u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m2 z a vdd vdd p w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
.ends
