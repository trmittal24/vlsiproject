* Tue Aug 10 11:21:07 CEST 2004
.subckt cgi2a_x2 a b c vdd vss z 
*SPICE circuit <cgi2a_x2> from XCircuit v3.10

m1 an a vss vss n w=30u l=2u ad='30u*5u+12p' as='30u*5u+12p' pd='30u*2+14u' ps='30u*2+14u'
m2 n3 b vss vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m3 an a vdd vdd p w=60u l=2u ad='60u*5u+12p' as='60u*5u+12p' pd='60u*2+14u' ps='60u*2+14u'
m4 n1 b vdd vdd p w=74u l=2u ad='74u*5u+12p' as='74u*5u+12p' pd='74u*2+14u' ps='74u*2+14u'
m5 n4 an vss vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m6 z c n3 vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m7 z b n2 vdd p w=74u l=2u ad='74u*5u+12p' as='74u*5u+12p' pd='74u*2+14u' ps='74u*2+14u'
m8 n2 an vdd vdd p w=74u l=2u ad='74u*5u+12p' as='74u*5u+12p' pd='74u*2+14u' ps='74u*2+14u'
m9 z c n1 vdd p w=74u l=2u ad='74u*5u+12p' as='74u*5u+12p' pd='74u*2+14u' ps='74u*2+14u'
m10 n1 an vdd vdd p w=74u l=2u ad='74u*5u+12p' as='74u*5u+12p' pd='74u*2+14u' ps='74u*2+14u'
m11 n3 an vss vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
.ends
