* Sun Apr  9 08:49:36 CEST 2006
.subckt oai21v0x4 a1 a2 b vdd vss z 
*SPICE circuit <oai21v0x4> from XCircuit v3.20

m1 n2 a1 vdd vdd p w=104u l=2u ad='104u*5u+12p' as='104u*5u+12p' pd='104u*2+14u' ps='104u*2+14u'
m2 z b vdd vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m3 n1 a2 vss vss n w=46u l=2u ad='46u*5u+12p' as='46u*5u+12p' pd='46u*2+14u' ps='46u*2+14u'
m4 n1 a1 vss vss n w=46u l=2u ad='46u*5u+12p' as='46u*5u+12p' pd='46u*2+14u' ps='46u*2+14u'
m5 z b n1 vss n w=49u l=2u ad='49u*5u+12p' as='49u*5u+12p' pd='49u*2+14u' ps='49u*2+14u'
m6 z a2 n2 vdd p w=104u l=2u ad='104u*5u+12p' as='104u*5u+12p' pd='104u*2+14u' ps='104u*2+14u'
.ends
