* Tue Dec 13 18:21:38 CET 2005
.subckt an2v0x4 a b vdd vss z 
*SPICE circuit <an2v0x4> from XCircuit v3.20

m1 z zn vdd vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m2 z zn vss vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m3 n1 a vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m4 zn a vdd vdd p w=25u l=2u ad='25u*5u+12p' as='25u*5u+12p' pd='25u*2+14u' ps='25u*2+14u'
m5 zn b n1 vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m6 zn b vdd vdd p w=25u l=2u ad='25u*5u+12p' as='25u*5u+12p' pd='25u*2+14u' ps='25u*2+14u'
.ends
