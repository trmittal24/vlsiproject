magic
tech scmos
timestamp 1521484183
use xnr2v8x05  xnr2v8x05_0
timestamp 1521484183
transform 1 0 4 0 1 4
box -4 -4 76 76
<< end >>
