* Spice description of nr3v1x05
* Spice driver version 134999461
* Date 17/05/2007 at  9:28:37
* vsclib 0.13um values
.subckt nr3v1x05 a b c vdd vss z
M01 vdd   a     n1    vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M02 vss   a     z     vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
M03 n1    b     05    vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M04 z     b     vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
M05 05    c     z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M06 vss   c     z     vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
C5  a     vss   0.475f
C3  b     vss   0.367f
C4  c     vss   0.369f
C2  z     vss   0.754f
.ends
