* Spice description of vfeed3
* Spice driver version 134999461
* Date 31/05/2007 at 21:36:00
* vxlib 0.13um values
.subckt vfeed3 vdd vss
.ends
