* Tue Dec 14 08:55:27 CET 2004
.subckt cgi2abv0x2 a b c vdd vss z 
*SPICE circuit <cgi2abv0x2> from XCircuit v3.20

m1 an a vss vss n w=22u l=2.3636u ad='22u*5u+12p' as='22u*5u+12p' pd='22u*2+14u' ps='22u*2+14u'
m2 bn b vss vss n w=22u l=2.3636u ad='22u*5u+12p' as='22u*5u+12p' pd='22u*2+14u' ps='22u*2+14u'
m3 an a vdd vdd p w=44u l=2.3636u ad='44u*5u+12p' as='44u*5u+12p' pd='44u*2+14u' ps='44u*2+14u'
m4 n3 bn vss vss n w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m5 bn b vdd vdd p w=44u l=2.3636u ad='44u*5u+12p' as='44u*5u+12p' pd='44u*2+14u' ps='44u*2+14u'
m6 n1 bn vdd vdd p w=54u l=2.3636u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m7 n2 an vdd vdd p w=54u l=2.3636u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m8 z bn n2 vdd p w=54u l=2.3636u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m9 n4 an vss vss n w=24u l=2.3636u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m10 z bn n4 vss n w=24u l=2.3636u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m11 z c n1 vdd p w=54u l=2.3636u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m12 n1 an vdd vdd p w=54u l=2.3636u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m13 n3 an vss vss n w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m14 z c n3 vss n w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
.ends
