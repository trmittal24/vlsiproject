* Tue Feb 20 08:57:11 CET 2007
.subckt xnr2v0x1 a b vdd vss z
*SPICE circuit <xnr2v0x1> from XCircuit v3.4 rev 26

m1 n1 an vdd vdd p w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m2 z b an vdd p w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m3 bn b vss vss n w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m4 an a vss vss n w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m5 z an bn vss n w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m6 an a vdd vdd p w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m7 bn b vdd vdd p w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m8 z bn an vss n w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m9 z bn n1 vdd p w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
.ends
