* Tue Aug 10 11:21:07 CEST 2004
.subckt nr3_x1 a b c vdd vss z 
*SPICE circuit <nr3_x1> from XCircuit v3.10

m1 z a vss vss n w=15u l=2.3636u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m2 z b vss vss n w=15u l=2.3636u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m3 z c vss vss n w=15u l=2.3636u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m4 z c n2 vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
m5 n2 b n1 vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
m6 n1 a vdd vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
.ends
