* SPICE3 file created from subcomp.ext - technology: scmos
.include t14y_tsmc_025_level3.txt

M1000 mux_0_vdd mux_0_mxn2v0x1_2_zn mux_0_o2 mux_0_mxn2v0x1_1_w_n4_32# pfet w=18u l=2u
+  ad=32118p pd=11574u as=102p ps=50u
M1001 mux_0_mxn2v0x1_2_a_21_50# mux_0_a2 mux_0_vdd mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1002 mux_0_mxn2v0x1_2_zn mux_0_s mux_0_mxn2v0x1_2_a_21_50# mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1003 mux_0_mxn2v0x1_2_a_38_50# mux_0_mxn2v0x1_2_sn mux_0_mxn2v0x1_2_zn mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1004 mux_0_vdd mux_0_b2 mux_0_mxn2v0x1_2_a_38_50# mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1005 mux_0_mxn2v0x1_2_sn mux_0_s mux_0_vdd mux_0_mxn2v0x1_1_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1006 mux_0_gnd mux_0_mxn2v0x1_2_zn mux_0_o2 mux_0_mxn2v0x1_2_w_n4_n4# nfet w=9u l=2u
+  ad=21409p pd=7648u as=57p ps=32u
M1007 mux_0_mxn2v0x1_2_a_21_12# mux_0_a2 mux_0_gnd mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1008 mux_0_mxn2v0x1_2_zn mux_0_mxn2v0x1_2_sn mux_0_mxn2v0x1_2_a_21_12# mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1009 mux_0_mxn2v0x1_2_a_38_12# mux_0_s mux_0_mxn2v0x1_2_zn mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1010 mux_0_gnd mux_0_b2 mux_0_mxn2v0x1_2_a_38_12# mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1011 mux_0_mxn2v0x1_2_sn mux_0_s mux_0_gnd mux_0_mxn2v0x1_2_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1012 mux_0_vdd mux_0_mxn2v0x1_1_zn mux_0_o1 mux_0_mxn2v0x1_1_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1013 mux_0_mxn2v0x1_1_a_21_50# mux_0_a1 mux_0_vdd mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1014 mux_0_mxn2v0x1_1_zn mux_0_s mux_0_mxn2v0x1_1_a_21_50# mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1015 mux_0_mxn2v0x1_1_a_38_50# mux_0_mxn2v0x1_1_sn mux_0_mxn2v0x1_1_zn mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1016 mux_0_vdd mux_0_b1 mux_0_mxn2v0x1_1_a_38_50# mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1017 mux_0_mxn2v0x1_1_sn mux_0_s mux_0_vdd mux_0_mxn2v0x1_1_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1018 mux_0_gnd mux_0_mxn2v0x1_1_zn mux_0_o1 mux_0_mxn2v0x1_0_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1019 mux_0_mxn2v0x1_1_a_21_12# mux_0_a1 mux_0_gnd mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1020 mux_0_mxn2v0x1_1_zn mux_0_mxn2v0x1_1_sn mux_0_mxn2v0x1_1_a_21_12# mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1021 mux_0_mxn2v0x1_1_a_38_12# mux_0_s mux_0_mxn2v0x1_1_zn mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1022 mux_0_gnd mux_0_b1 mux_0_mxn2v0x1_1_a_38_12# mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1023 mux_0_mxn2v0x1_1_sn mux_0_s mux_0_gnd mux_0_mxn2v0x1_0_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1024 mux_0_vdd mux_0_mxn2v0x1_0_zn mux_0_o0 mux_0_mxn2v0x1_0_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1025 mux_0_mxn2v0x1_0_a_21_50# mux_0_a0 mux_0_vdd mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1026 mux_0_mxn2v0x1_0_zn mux_0_s mux_0_mxn2v0x1_0_a_21_50# mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1027 mux_0_mxn2v0x1_0_a_38_50# mux_0_mxn2v0x1_0_sn mux_0_mxn2v0x1_0_zn mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1028 mux_0_vdd mux_0_b0 mux_0_mxn2v0x1_0_a_38_50# mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1029 mux_0_mxn2v0x1_0_sn mux_0_s mux_0_vdd mux_0_mxn2v0x1_0_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1030 mux_0_gnd mux_0_mxn2v0x1_0_zn mux_0_o0 mux_0_mxn2v0x1_0_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1031 mux_0_mxn2v0x1_0_a_21_12# mux_0_a0 mux_0_gnd mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1032 mux_0_mxn2v0x1_0_zn mux_0_mxn2v0x1_0_sn mux_0_mxn2v0x1_0_a_21_12# mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1033 mux_0_mxn2v0x1_0_a_38_12# mux_0_s mux_0_mxn2v0x1_0_zn mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1034 mux_0_gnd mux_0_b0 mux_0_mxn2v0x1_0_a_38_12# mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1035 mux_0_mxn2v0x1_0_sn mux_0_s mux_0_gnd mux_0_mxn2v0x1_0_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1036 mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_2_zn mux_0_a2 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1037 totdiff3_0_mux_0_mxn2v0x1_2_a_21_50# totdiff3_0_mux_0_a2 mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1038 totdiff3_0_mux_0_mxn2v0x1_2_zn totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_2_a_21_50# totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1039 totdiff3_0_mux_0_mxn2v0x1_2_a_38_50# totdiff3_0_mux_0_mxn2v0x1_2_sn totdiff3_0_mux_0_mxn2v0x1_2_zn totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1040 mux_0_vdd totdiff3_0_mux_0_b2 totdiff3_0_mux_0_mxn2v0x1_2_a_38_50# totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1041 totdiff3_0_mux_0_mxn2v0x1_2_sn totdiff3_0_mux_0_s mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1042 mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_2_zn mux_0_a2 totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1043 totdiff3_0_mux_0_mxn2v0x1_2_a_21_12# totdiff3_0_mux_0_a2 mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1044 totdiff3_0_mux_0_mxn2v0x1_2_zn totdiff3_0_mux_0_mxn2v0x1_2_sn totdiff3_0_mux_0_mxn2v0x1_2_a_21_12# totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1045 totdiff3_0_mux_0_mxn2v0x1_2_a_38_12# totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_2_zn totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1046 mux_0_gnd totdiff3_0_mux_0_b2 totdiff3_0_mux_0_mxn2v0x1_2_a_38_12# totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1047 totdiff3_0_mux_0_mxn2v0x1_2_sn totdiff3_0_mux_0_s mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1048 mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_1_zn mux_0_a1 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1049 totdiff3_0_mux_0_mxn2v0x1_1_a_21_50# totdiff3_0_mux_0_a1 mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1050 totdiff3_0_mux_0_mxn2v0x1_1_zn totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_1_a_21_50# totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1051 totdiff3_0_mux_0_mxn2v0x1_1_a_38_50# totdiff3_0_mux_0_mxn2v0x1_1_sn totdiff3_0_mux_0_mxn2v0x1_1_zn totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1052 mux_0_vdd totdiff3_0_mux_0_b1 totdiff3_0_mux_0_mxn2v0x1_1_a_38_50# totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1053 totdiff3_0_mux_0_mxn2v0x1_1_sn totdiff3_0_mux_0_s mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1054 mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_1_zn mux_0_a1 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1055 totdiff3_0_mux_0_mxn2v0x1_1_a_21_12# totdiff3_0_mux_0_a1 mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1056 totdiff3_0_mux_0_mxn2v0x1_1_zn totdiff3_0_mux_0_mxn2v0x1_1_sn totdiff3_0_mux_0_mxn2v0x1_1_a_21_12# totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1057 totdiff3_0_mux_0_mxn2v0x1_1_a_38_12# totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_1_zn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1058 mux_0_gnd totdiff3_0_mux_0_b1 totdiff3_0_mux_0_mxn2v0x1_1_a_38_12# totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1059 totdiff3_0_mux_0_mxn2v0x1_1_sn totdiff3_0_mux_0_s mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1060 mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_0_zn mux_0_a0 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1061 totdiff3_0_mux_0_mxn2v0x1_0_a_21_50# totdiff3_0_mux_0_a0 mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1062 totdiff3_0_mux_0_mxn2v0x1_0_zn totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_0_a_21_50# totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1063 totdiff3_0_mux_0_mxn2v0x1_0_a_38_50# totdiff3_0_mux_0_mxn2v0x1_0_sn totdiff3_0_mux_0_mxn2v0x1_0_zn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1064 mux_0_vdd totdiff3_0_mux_0_b0 totdiff3_0_mux_0_mxn2v0x1_0_a_38_50# totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1065 totdiff3_0_mux_0_mxn2v0x1_0_sn totdiff3_0_mux_0_s mux_0_vdd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1066 mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_0_zn mux_0_a0 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1067 totdiff3_0_mux_0_mxn2v0x1_0_a_21_12# totdiff3_0_mux_0_a0 mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1068 totdiff3_0_mux_0_mxn2v0x1_0_zn totdiff3_0_mux_0_mxn2v0x1_0_sn totdiff3_0_mux_0_mxn2v0x1_0_a_21_12# totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1069 totdiff3_0_mux_0_mxn2v0x1_0_a_38_12# totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_0_zn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1070 mux_0_gnd totdiff3_0_mux_0_b0 totdiff3_0_mux_0_mxn2v0x1_0_a_38_12# totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1071 totdiff3_0_mux_0_mxn2v0x1_0_sn totdiff3_0_mux_0_s mux_0_gnd totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1072 mux_0_vdd totdiff3_0_diff2_2_an2v0x2_2_zn totdiff3_0_diff2_2_an2v0x2_2_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1073 totdiff3_0_diff2_2_an2v0x2_2_zn totdiff3_0_diff2_2_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1074 mux_0_vdd totdiff3_0_diff2_2_in_2c totdiff3_0_diff2_2_an2v0x2_2_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1075 mux_0_gnd totdiff3_0_diff2_2_an2v0x2_2_zn totdiff3_0_diff2_2_an2v0x2_2_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1076 totdiff3_0_diff2_2_an2v0x2_2_a_24_13# totdiff3_0_diff2_2_an2v0x2_2_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1077 totdiff3_0_diff2_2_an2v0x2_2_zn totdiff3_0_diff2_2_in_2c totdiff3_0_diff2_2_an2v0x2_2_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1078 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_mux_0_b2 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1079 totdiff3_0_mux_0_b2 totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_diff2_2_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1080 totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_b2 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1081 totdiff3_0_mux_0_b2 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_diff2_2_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1082 totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_diff2_2_in_2c mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1083 mux_0_vdd totdiff3_0_diff2_2_in_2c totdiff3_0_diff2_2_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1084 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_diff2_2_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1085 mux_0_vdd totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_diff2_2_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1086 totdiff3_0_diff2_2_xor2v2x2_0_a_13_13# totdiff3_0_diff2_2_xor2v2x2_0_an mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1087 totdiff3_0_mux_0_b2 totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_diff2_2_xor2v2x2_0_a_13_13# mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1088 totdiff3_0_diff2_2_xor2v2x2_0_a_30_13# totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_mux_0_b2 mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1089 mux_0_gnd totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_diff2_2_xor2v2x2_0_a_30_13# mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1090 totdiff3_0_diff2_2_xor2v2x2_0_bn totdiff3_0_diff2_2_in_2c mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1091 totdiff3_0_mux_0_b2 totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_diff2_2_xor2v2x2_0_bn mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1092 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_diff2_2_in_2c totdiff3_0_mux_0_b2 mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1093 mux_0_gnd totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_diff2_2_xor2v2x2_0_an mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1094 totdiff3_0_mux_0_s totdiff3_0_diff2_2_or2v0x3_0_zn mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1095 mux_0_vdd totdiff3_0_diff2_2_or2v0x3_0_zn totdiff3_0_mux_0_s mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1096 totdiff3_0_diff2_2_or2v0x3_0_a_31_39# totdiff3_0_diff2_2_an2v0x2_1_z mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1097 totdiff3_0_diff2_2_or2v0x3_0_zn totdiff3_0_diff2_2_an2v0x2_0_z totdiff3_0_diff2_2_or2v0x3_0_a_31_39# mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1098 totdiff3_0_diff2_2_or2v0x3_0_a_48_39# totdiff3_0_diff2_2_an2v0x2_0_z totdiff3_0_diff2_2_or2v0x3_0_zn mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1099 mux_0_vdd totdiff3_0_diff2_2_an2v0x2_1_z totdiff3_0_diff2_2_or2v0x3_0_a_48_39# mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1100 mux_0_gnd totdiff3_0_diff2_2_or2v0x3_0_zn totdiff3_0_mux_0_s mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1101 totdiff3_0_diff2_2_or2v0x3_0_zn totdiff3_0_diff2_2_an2v0x2_1_z mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1102 mux_0_gnd totdiff3_0_diff2_2_an2v0x2_0_z totdiff3_0_diff2_2_or2v0x3_0_zn mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1103 mux_0_vdd totdiff3_0_diff2_2_an2v0x2_1_zn totdiff3_0_diff2_2_an2v0x2_1_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1104 totdiff3_0_diff2_2_an2v0x2_1_zn totdiff3_0_diff2_2_an2v0x2_1_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1105 mux_0_vdd totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_an2v0x2_1_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1106 mux_0_gnd totdiff3_0_diff2_2_an2v0x2_1_zn totdiff3_0_diff2_2_an2v0x2_1_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1107 totdiff3_0_diff2_2_an2v0x2_1_a_24_13# totdiff3_0_diff2_2_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1108 totdiff3_0_diff2_2_an2v0x2_1_zn totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_an2v0x2_1_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1109 mux_0_vdd totdiff3_0_diff2_2_an2v0x2_0_zn totdiff3_0_diff2_2_an2v0x2_0_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1110 totdiff3_0_diff2_2_an2v0x2_0_zn totdiff3_0_diff2_2_in_c mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1111 mux_0_vdd totdiff3_0_diff2_2_an2v0x2_0_b totdiff3_0_diff2_2_an2v0x2_0_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1112 mux_0_gnd totdiff3_0_diff2_2_an2v0x2_0_zn totdiff3_0_diff2_2_an2v0x2_0_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1113 totdiff3_0_diff2_2_an2v0x2_0_a_24_13# totdiff3_0_diff2_2_in_c mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1114 totdiff3_0_diff2_2_an2v0x2_0_zn totdiff3_0_diff2_2_an2v0x2_0_b totdiff3_0_diff2_2_an2v0x2_0_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1115 mux_0_vdd totdiff3_0_diff2_2_xnr2v8x05_0_zn totdiff3_0_diff2_2_an2v0x2_0_b mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1116 totdiff3_0_diff2_2_xnr2v8x05_0_an totdiff3_0_diff2_2_in_a mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1117 totdiff3_0_diff2_2_xnr2v8x05_0_zn totdiff3_0_diff2_2_xnr2v8x05_0_bn totdiff3_0_diff2_2_xnr2v8x05_0_an mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1118 totdiff3_0_diff2_2_xnr2v8x05_0_ai totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_xnr2v8x05_0_zn mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1119 mux_0_vdd totdiff3_0_diff2_2_xnr2v8x05_0_an totdiff3_0_diff2_2_xnr2v8x05_0_ai mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1120 totdiff3_0_diff2_2_xnr2v8x05_0_bn totdiff3_0_diff2_2_in_b mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1121 mux_0_gnd totdiff3_0_diff2_2_xnr2v8x05_0_zn totdiff3_0_diff2_2_an2v0x2_0_b mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1122 totdiff3_0_diff2_2_xnr2v8x05_0_an totdiff3_0_diff2_2_in_a mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1123 totdiff3_0_diff2_2_xnr2v8x05_0_zn totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_xnr2v8x05_0_an mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1124 totdiff3_0_diff2_2_xnr2v8x05_0_ai totdiff3_0_diff2_2_xnr2v8x05_0_bn totdiff3_0_diff2_2_xnr2v8x05_0_zn mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1125 mux_0_gnd totdiff3_0_diff2_2_xnr2v8x05_0_an totdiff3_0_diff2_2_xnr2v8x05_0_ai mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1126 totdiff3_0_diff2_2_xnr2v8x05_0_bn totdiff3_0_diff2_2_in_b mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1127 totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_a2 mux_0_vdd mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1128 mux_0_vdd totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_an2v0x2_2_a mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1129 totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_mux_0_a2 mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1130 mux_0_gnd totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_an2v0x2_2_a mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1131 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_a2 mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1132 totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_xor3v1x2_0_cn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1133 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_mux_0_a2 mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1134 totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_xor3v1x2_0_zn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1135 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_in_c mux_0_vdd mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1136 mux_0_vdd totdiff3_0_diff2_2_in_c totdiff3_0_diff2_2_xor3v1x2_0_cn mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1137 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_xor3v1x2_0_iz mux_0_vdd mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1138 mux_0_vdd totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_diff2_2_xor3v1x2_0_zn mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1139 totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_diff2_2_an2v0x2_1_a totdiff3_0_diff2_2_xor3v1x2_0_bn mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1140 totdiff3_0_diff2_2_an2v0x2_1_a totdiff3_0_diff2_2_xor3v1x2_0_bn totdiff3_0_diff2_2_xor3v1x2_0_iz mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1141 mux_0_vdd totdiff3_0_diff2_2_in_a totdiff3_0_diff2_2_an2v0x2_1_a mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1142 totdiff3_0_diff2_2_xor3v1x2_0_bn totdiff3_0_diff2_2_in_b mux_0_vdd mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1143 mux_0_vdd totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_xor3v1x2_0_bn mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1144 totdiff3_0_diff2_2_xor3v1x2_0_a_11_12# totdiff3_0_diff2_2_xor3v1x2_0_cn mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1145 totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_xor3v1x2_0_a_11_12# mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1146 totdiff3_0_diff2_2_xor3v1x2_0_a_28_12# totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_a2 mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1147 mux_0_gnd totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_xor3v1x2_0_a_28_12# mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1148 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_xor3v1x2_0_iz mux_0_gnd mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1149 totdiff3_0_mux_0_a2 totdiff3_0_diff2_2_in_c totdiff3_0_diff2_2_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1150 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_in_c totdiff3_0_mux_0_a2 mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1151 mux_0_gnd totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_diff2_2_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1152 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_in_c mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1153 mux_0_gnd totdiff3_0_diff2_2_in_c totdiff3_0_diff2_2_xor3v1x2_0_cn mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1154 totdiff3_0_diff2_2_xor3v1x2_0_a_115_7# totdiff3_0_diff2_2_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1155 totdiff3_0_diff2_2_xor3v1x2_0_iz totdiff3_0_diff2_2_xor3v1x2_0_bn totdiff3_0_diff2_2_xor3v1x2_0_a_115_7# mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1156 totdiff3_0_diff2_2_an2v0x2_1_a totdiff3_0_diff2_2_in_b totdiff3_0_diff2_2_xor3v1x2_0_iz mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1157 mux_0_gnd totdiff3_0_diff2_2_in_a totdiff3_0_diff2_2_an2v0x2_1_a mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1158 totdiff3_0_diff2_2_xor3v1x2_0_bn totdiff3_0_diff2_2_in_b mux_0_gnd mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1159 mux_0_vdd totdiff3_0_diff2_1_an2v0x2_2_zn totdiff3_0_diff2_2_in_2c mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1160 totdiff3_0_diff2_1_an2v0x2_2_zn totdiff3_0_diff2_1_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1161 mux_0_vdd totdiff3_0_diff2_1_in_2c totdiff3_0_diff2_1_an2v0x2_2_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1162 mux_0_gnd totdiff3_0_diff2_1_an2v0x2_2_zn totdiff3_0_diff2_2_in_2c mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1163 totdiff3_0_diff2_1_an2v0x2_2_a_24_13# totdiff3_0_diff2_1_an2v0x2_2_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1164 totdiff3_0_diff2_1_an2v0x2_2_zn totdiff3_0_diff2_1_in_2c totdiff3_0_diff2_1_an2v0x2_2_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1165 totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_mux_0_b1 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1166 totdiff3_0_mux_0_b1 totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_diff2_1_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1167 totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_mux_0_b1 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1168 totdiff3_0_mux_0_b1 totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_diff2_1_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1169 totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_diff2_1_in_2c mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1170 mux_0_vdd totdiff3_0_diff2_1_in_2c totdiff3_0_diff2_1_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1171 totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_diff2_1_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1172 mux_0_vdd totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_diff2_1_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1173 totdiff3_0_diff2_1_xor2v2x2_0_a_13_13# totdiff3_0_diff2_1_xor2v2x2_0_an mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1174 totdiff3_0_mux_0_b1 totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_diff2_1_xor2v2x2_0_a_13_13# mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1175 totdiff3_0_diff2_1_xor2v2x2_0_a_30_13# totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_mux_0_b1 mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1176 mux_0_gnd totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_diff2_1_xor2v2x2_0_a_30_13# mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1177 totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_diff2_1_in_2c mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1178 totdiff3_0_mux_0_b1 totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_diff2_1_xor2v2x2_0_bn mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1179 totdiff3_0_diff2_1_xor2v2x2_0_an totdiff3_0_diff2_1_in_2c totdiff3_0_mux_0_b1 mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1180 mux_0_gnd totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_diff2_1_xor2v2x2_0_an mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1181 totdiff3_0_diff2_2_in_c totdiff3_0_diff2_1_or2v0x3_0_zn mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1182 mux_0_vdd totdiff3_0_diff2_1_or2v0x3_0_zn totdiff3_0_diff2_2_in_c mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1183 totdiff3_0_diff2_1_or2v0x3_0_a_31_39# totdiff3_0_diff2_1_an2v0x2_1_z mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1184 totdiff3_0_diff2_1_or2v0x3_0_zn totdiff3_0_diff2_1_an2v0x2_0_z totdiff3_0_diff2_1_or2v0x3_0_a_31_39# mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1185 totdiff3_0_diff2_1_or2v0x3_0_a_48_39# totdiff3_0_diff2_1_an2v0x2_0_z totdiff3_0_diff2_1_or2v0x3_0_zn mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1186 mux_0_vdd totdiff3_0_diff2_1_an2v0x2_1_z totdiff3_0_diff2_1_or2v0x3_0_a_48_39# mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1187 mux_0_gnd totdiff3_0_diff2_1_or2v0x3_0_zn totdiff3_0_diff2_2_in_c mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1188 totdiff3_0_diff2_1_or2v0x3_0_zn totdiff3_0_diff2_1_an2v0x2_1_z mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1189 mux_0_gnd totdiff3_0_diff2_1_an2v0x2_0_z totdiff3_0_diff2_1_or2v0x3_0_zn mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1190 mux_0_vdd totdiff3_0_diff2_1_an2v0x2_1_zn totdiff3_0_diff2_1_an2v0x2_1_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1191 totdiff3_0_diff2_1_an2v0x2_1_zn totdiff3_0_diff2_1_an2v0x2_1_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1192 mux_0_vdd totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_an2v0x2_1_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1193 mux_0_gnd totdiff3_0_diff2_1_an2v0x2_1_zn totdiff3_0_diff2_1_an2v0x2_1_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1194 totdiff3_0_diff2_1_an2v0x2_1_a_24_13# totdiff3_0_diff2_1_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1195 totdiff3_0_diff2_1_an2v0x2_1_zn totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_an2v0x2_1_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1196 mux_0_vdd totdiff3_0_diff2_1_an2v0x2_0_zn totdiff3_0_diff2_1_an2v0x2_0_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1197 totdiff3_0_diff2_1_an2v0x2_0_zn totdiff3_0_diff2_1_in_c mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1198 mux_0_vdd totdiff3_0_diff2_1_an2v0x2_0_b totdiff3_0_diff2_1_an2v0x2_0_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1199 mux_0_gnd totdiff3_0_diff2_1_an2v0x2_0_zn totdiff3_0_diff2_1_an2v0x2_0_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1200 totdiff3_0_diff2_1_an2v0x2_0_a_24_13# totdiff3_0_diff2_1_in_c mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1201 totdiff3_0_diff2_1_an2v0x2_0_zn totdiff3_0_diff2_1_an2v0x2_0_b totdiff3_0_diff2_1_an2v0x2_0_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1202 mux_0_vdd totdiff3_0_diff2_1_xnr2v8x05_0_zn totdiff3_0_diff2_1_an2v0x2_0_b mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1203 totdiff3_0_diff2_1_xnr2v8x05_0_an totdiff3_0_diff2_1_in_a mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1204 totdiff3_0_diff2_1_xnr2v8x05_0_zn totdiff3_0_diff2_1_xnr2v8x05_0_bn totdiff3_0_diff2_1_xnr2v8x05_0_an mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1205 totdiff3_0_diff2_1_xnr2v8x05_0_ai totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_xnr2v8x05_0_zn mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1206 mux_0_vdd totdiff3_0_diff2_1_xnr2v8x05_0_an totdiff3_0_diff2_1_xnr2v8x05_0_ai mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1207 totdiff3_0_diff2_1_xnr2v8x05_0_bn totdiff3_0_diff2_1_in_b mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1208 mux_0_gnd totdiff3_0_diff2_1_xnr2v8x05_0_zn totdiff3_0_diff2_1_an2v0x2_0_b mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1209 totdiff3_0_diff2_1_xnr2v8x05_0_an totdiff3_0_diff2_1_in_a mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1210 totdiff3_0_diff2_1_xnr2v8x05_0_zn totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_xnr2v8x05_0_an mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1211 totdiff3_0_diff2_1_xnr2v8x05_0_ai totdiff3_0_diff2_1_xnr2v8x05_0_bn totdiff3_0_diff2_1_xnr2v8x05_0_zn mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1212 mux_0_gnd totdiff3_0_diff2_1_xnr2v8x05_0_an totdiff3_0_diff2_1_xnr2v8x05_0_ai mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1213 totdiff3_0_diff2_1_xnr2v8x05_0_bn totdiff3_0_diff2_1_in_b mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1214 totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_a1 mux_0_vdd mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1215 mux_0_vdd totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_an2v0x2_2_a mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1216 totdiff3_0_diff2_1_an2v0x2_2_a totdiff3_0_mux_0_a1 mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1217 mux_0_gnd totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_an2v0x2_2_a mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1218 totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_a1 mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1219 totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_xor3v1x2_0_cn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1220 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_mux_0_a1 mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1221 totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_diff2_1_xor3v1x2_0_zn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1222 totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_diff2_1_in_c mux_0_vdd mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1223 mux_0_vdd totdiff3_0_diff2_1_in_c totdiff3_0_diff2_1_xor3v1x2_0_cn mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1224 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_xor3v1x2_0_iz mux_0_vdd mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1225 mux_0_vdd totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_diff2_1_xor3v1x2_0_zn mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1226 totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_diff2_1_an2v0x2_1_a totdiff3_0_diff2_1_xor3v1x2_0_bn mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1227 totdiff3_0_diff2_1_an2v0x2_1_a totdiff3_0_diff2_1_xor3v1x2_0_bn totdiff3_0_diff2_1_xor3v1x2_0_iz mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1228 mux_0_vdd totdiff3_0_diff2_1_in_a totdiff3_0_diff2_1_an2v0x2_1_a mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1229 totdiff3_0_diff2_1_xor3v1x2_0_bn totdiff3_0_diff2_1_in_b mux_0_vdd mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1230 mux_0_vdd totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_xor3v1x2_0_bn mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1231 totdiff3_0_diff2_1_xor3v1x2_0_a_11_12# totdiff3_0_diff2_1_xor3v1x2_0_cn mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1232 totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_xor3v1x2_0_a_11_12# mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1233 totdiff3_0_diff2_1_xor3v1x2_0_a_28_12# totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_a1 mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1234 mux_0_gnd totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_diff2_1_xor3v1x2_0_a_28_12# mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1235 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_xor3v1x2_0_iz mux_0_gnd mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1236 totdiff3_0_mux_0_a1 totdiff3_0_diff2_1_in_c totdiff3_0_diff2_1_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1237 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_in_c totdiff3_0_mux_0_a1 mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1238 mux_0_gnd totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_diff2_1_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1239 totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_diff2_1_in_c mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1240 mux_0_gnd totdiff3_0_diff2_1_in_c totdiff3_0_diff2_1_xor3v1x2_0_cn mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1241 totdiff3_0_diff2_1_xor3v1x2_0_a_115_7# totdiff3_0_diff2_1_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1242 totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_diff2_1_xor3v1x2_0_bn totdiff3_0_diff2_1_xor3v1x2_0_a_115_7# mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1243 totdiff3_0_diff2_1_an2v0x2_1_a totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_xor3v1x2_0_iz mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1244 mux_0_gnd totdiff3_0_diff2_1_in_a totdiff3_0_diff2_1_an2v0x2_1_a mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1245 totdiff3_0_diff2_1_xor3v1x2_0_bn totdiff3_0_diff2_1_in_b mux_0_gnd mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1246 mux_0_vdd totdiff3_0_diff2_0_an2v0x2_2_zn totdiff3_0_diff2_1_in_2c mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1247 totdiff3_0_diff2_0_an2v0x2_2_zn totdiff3_0_diff2_0_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1248 mux_0_vdd mux_0_vdd totdiff3_0_diff2_0_an2v0x2_2_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1249 mux_0_gnd totdiff3_0_diff2_0_an2v0x2_2_zn totdiff3_0_diff2_1_in_2c mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1250 totdiff3_0_diff2_0_an2v0x2_2_a_24_13# totdiff3_0_diff2_0_an2v0x2_2_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1251 totdiff3_0_diff2_0_an2v0x2_2_zn mux_0_vdd totdiff3_0_diff2_0_an2v0x2_2_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1252 totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_b0 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1253 totdiff3_0_mux_0_b0 totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_diff2_0_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1254 totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_mux_0_b0 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1255 totdiff3_0_mux_0_b0 totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_diff2_0_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1256 totdiff3_0_diff2_0_xor2v2x2_0_bn mux_0_vdd mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1257 mux_0_vdd mux_0_vdd totdiff3_0_diff2_0_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1258 totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_diff2_0_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1259 mux_0_vdd totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_diff2_0_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1260 totdiff3_0_diff2_0_xor2v2x2_0_a_13_13# totdiff3_0_diff2_0_xor2v2x2_0_an mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1261 totdiff3_0_mux_0_b0 totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_diff2_0_xor2v2x2_0_a_13_13# mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1262 totdiff3_0_diff2_0_xor2v2x2_0_a_30_13# totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_mux_0_b0 mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1263 mux_0_gnd totdiff3_0_diff2_0_xor2v2x2_0_an totdiff3_0_diff2_0_xor2v2x2_0_a_30_13# mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1264 totdiff3_0_diff2_0_xor2v2x2_0_bn mux_0_vdd mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1265 totdiff3_0_mux_0_b0 totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_diff2_0_xor2v2x2_0_bn mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1266 totdiff3_0_diff2_0_xor2v2x2_0_an mux_0_vdd totdiff3_0_mux_0_b0 mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1267 mux_0_gnd totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_diff2_0_xor2v2x2_0_an mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1268 totdiff3_0_diff2_1_in_c totdiff3_0_diff2_0_or2v0x3_0_zn mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1269 mux_0_vdd totdiff3_0_diff2_0_or2v0x3_0_zn totdiff3_0_diff2_1_in_c mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1270 totdiff3_0_diff2_0_or2v0x3_0_a_31_39# totdiff3_0_diff2_0_an2v0x2_1_z mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1271 totdiff3_0_diff2_0_or2v0x3_0_zn totdiff3_0_diff2_0_an2v0x2_0_z totdiff3_0_diff2_0_or2v0x3_0_a_31_39# mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1272 totdiff3_0_diff2_0_or2v0x3_0_a_48_39# totdiff3_0_diff2_0_an2v0x2_0_z totdiff3_0_diff2_0_or2v0x3_0_zn mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1273 mux_0_vdd totdiff3_0_diff2_0_an2v0x2_1_z totdiff3_0_diff2_0_or2v0x3_0_a_48_39# mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1274 mux_0_gnd totdiff3_0_diff2_0_or2v0x3_0_zn totdiff3_0_diff2_1_in_c mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1275 totdiff3_0_diff2_0_or2v0x3_0_zn totdiff3_0_diff2_0_an2v0x2_1_z mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1276 mux_0_gnd totdiff3_0_diff2_0_an2v0x2_0_z totdiff3_0_diff2_0_or2v0x3_0_zn mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1277 mux_0_vdd totdiff3_0_diff2_0_an2v0x2_1_zn totdiff3_0_diff2_0_an2v0x2_1_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1278 totdiff3_0_diff2_0_an2v0x2_1_zn totdiff3_0_diff2_0_an2v0x2_1_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1279 mux_0_vdd totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_an2v0x2_1_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1280 mux_0_gnd totdiff3_0_diff2_0_an2v0x2_1_zn totdiff3_0_diff2_0_an2v0x2_1_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1281 totdiff3_0_diff2_0_an2v0x2_1_a_24_13# totdiff3_0_diff2_0_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1282 totdiff3_0_diff2_0_an2v0x2_1_zn totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_an2v0x2_1_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1283 mux_0_vdd totdiff3_0_diff2_0_an2v0x2_0_zn totdiff3_0_diff2_0_an2v0x2_0_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1284 totdiff3_0_diff2_0_an2v0x2_0_zn mux_0_gnd mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1285 mux_0_vdd totdiff3_0_diff2_0_an2v0x2_0_b totdiff3_0_diff2_0_an2v0x2_0_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1286 mux_0_gnd totdiff3_0_diff2_0_an2v0x2_0_zn totdiff3_0_diff2_0_an2v0x2_0_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1287 totdiff3_0_diff2_0_an2v0x2_0_a_24_13# mux_0_gnd mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1288 totdiff3_0_diff2_0_an2v0x2_0_zn totdiff3_0_diff2_0_an2v0x2_0_b totdiff3_0_diff2_0_an2v0x2_0_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1289 mux_0_vdd totdiff3_0_diff2_0_xnr2v8x05_0_zn totdiff3_0_diff2_0_an2v0x2_0_b mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1290 totdiff3_0_diff2_0_xnr2v8x05_0_an totdiff3_0_diff2_0_in_a mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1291 totdiff3_0_diff2_0_xnr2v8x05_0_zn totdiff3_0_diff2_0_xnr2v8x05_0_bn totdiff3_0_diff2_0_xnr2v8x05_0_an mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1292 totdiff3_0_diff2_0_xnr2v8x05_0_ai totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_xnr2v8x05_0_zn mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1293 mux_0_vdd totdiff3_0_diff2_0_xnr2v8x05_0_an totdiff3_0_diff2_0_xnr2v8x05_0_ai mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1294 totdiff3_0_diff2_0_xnr2v8x05_0_bn totdiff3_0_diff2_0_in_b mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1295 mux_0_gnd totdiff3_0_diff2_0_xnr2v8x05_0_zn totdiff3_0_diff2_0_an2v0x2_0_b mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1296 totdiff3_0_diff2_0_xnr2v8x05_0_an totdiff3_0_diff2_0_in_a mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1297 totdiff3_0_diff2_0_xnr2v8x05_0_zn totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_xnr2v8x05_0_an mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1298 totdiff3_0_diff2_0_xnr2v8x05_0_ai totdiff3_0_diff2_0_xnr2v8x05_0_bn totdiff3_0_diff2_0_xnr2v8x05_0_zn mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1299 mux_0_gnd totdiff3_0_diff2_0_xnr2v8x05_0_an totdiff3_0_diff2_0_xnr2v8x05_0_ai mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1300 totdiff3_0_diff2_0_xnr2v8x05_0_bn totdiff3_0_diff2_0_in_b mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1301 totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_a0 mux_0_vdd mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1302 mux_0_vdd totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_an2v0x2_2_a mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1303 totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_mux_0_a0 mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1304 mux_0_gnd totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_an2v0x2_2_a mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1305 totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_a0 mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1306 totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_diff2_0_xor3v1x2_0_cn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1307 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_mux_0_a0 mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1308 totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_diff2_0_xor3v1x2_0_zn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1309 totdiff3_0_diff2_0_xor3v1x2_0_cn mux_0_gnd mux_0_vdd mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1310 mux_0_vdd mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_cn mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1311 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_diff2_0_xor3v1x2_0_iz mux_0_vdd mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1312 mux_0_vdd totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_diff2_0_xor3v1x2_0_zn mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1313 totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_diff2_0_xor3v1x2_0_bn mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1314 totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_diff2_0_xor3v1x2_0_iz mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1315 mux_0_vdd totdiff3_0_diff2_0_in_a totdiff3_0_diff2_0_an2v0x2_1_a mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1316 totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_diff2_0_in_b mux_0_vdd mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1317 mux_0_vdd totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_xor3v1x2_0_bn mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1318 totdiff3_0_diff2_0_xor3v1x2_0_a_11_12# totdiff3_0_diff2_0_xor3v1x2_0_cn mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1319 totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_diff2_0_xor3v1x2_0_a_11_12# mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1320 totdiff3_0_diff2_0_xor3v1x2_0_a_28_12# totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_mux_0_a0 mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1321 mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_diff2_0_xor3v1x2_0_a_28_12# mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1322 totdiff3_0_diff2_0_xor3v1x2_0_zn totdiff3_0_diff2_0_xor3v1x2_0_iz mux_0_gnd mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1323 totdiff3_0_mux_0_a0 mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1324 totdiff3_0_diff2_0_xor3v1x2_0_zn mux_0_gnd totdiff3_0_mux_0_a0 mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1325 mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_diff2_0_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1326 totdiff3_0_diff2_0_xor3v1x2_0_cn mux_0_gnd mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1327 mux_0_gnd mux_0_gnd totdiff3_0_diff2_0_xor3v1x2_0_cn mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1328 totdiff3_0_diff2_0_xor3v1x2_0_a_115_7# totdiff3_0_diff2_0_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1329 totdiff3_0_diff2_0_xor3v1x2_0_iz totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_diff2_0_xor3v1x2_0_a_115_7# mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1330 totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_xor3v1x2_0_iz mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1331 mux_0_gnd totdiff3_0_diff2_0_in_a totdiff3_0_diff2_0_an2v0x2_1_a mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1332 totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_diff2_0_in_b mux_0_gnd mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1333 comp_0_nd3v0x2_0_z comp_0_nr3v0x2_0_z mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=14u l=2u
+  ad=392p pd=120u as=0p ps=0u
M1334 mux_0_vdd comp_0_nr3v0x2_0_z comp_0_nd3v0x2_0_z comp_0_an3v0x2_2_w_n4_32# pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1335 comp_0_nd3v0x2_0_z comp_0_nd3v0x2_0_c mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1336 mux_0_vdd comp_0_nd3v0x2_0_a comp_0_nd3v0x2_0_z comp_0_an3v0x2_2_w_n4_32# pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1337 comp_0_nd3v0x2_0_a_14_12# comp_0_nd3v0x2_0_a mux_0_gnd mux_0_gnd nfet w=14u l=2u
+  ad=70p pd=38u as=0p ps=0u
M1338 comp_0_nd3v0x2_0_a_21_12# comp_0_nr3v0x2_0_z comp_0_nd3v0x2_0_a_14_12# mux_0_gnd nfet w=14u l=2u
+  ad=70p pd=38u as=0p ps=0u
M1339 comp_0_nd3v0x2_0_z comp_0_nd3v0x2_0_c comp_0_nd3v0x2_0_a_21_12# mux_0_gnd nfet w=14u l=2u
+  ad=112p pd=44u as=0p ps=0u
M1340 comp_0_nd3v0x2_0_a_38_12# comp_0_nd3v0x2_0_c comp_0_nd3v0x2_0_z mux_0_gnd nfet w=14u l=2u
+  ad=70p pd=38u as=0p ps=0u
M1341 comp_0_nd3v0x2_0_a_45_12# comp_0_nr3v0x2_0_z comp_0_nd3v0x2_0_a_38_12# mux_0_gnd nfet w=14u l=2u
+  ad=70p pd=38u as=0p ps=0u
M1342 mux_0_gnd comp_0_nd3v0x2_0_a comp_0_nd3v0x2_0_a_45_12# mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1343 mux_0_vdd comp_0_an3v0x2_1_zn comp_0_nr2v0x2_1_a comp_0_an3v0x2_2_w_n4_32# pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1344 comp_0_an3v0x2_1_zn comp_0_an3v0x2_1_a mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=17u l=2u
+  ad=233p pd=98u as=0p ps=0u
M1345 mux_0_vdd comp_0_an3v0x2_2_b comp_0_an3v0x2_1_zn comp_0_an3v0x2_2_w_n4_32# pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1346 comp_0_an3v0x2_1_zn mux_0_a2 mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1347 mux_0_gnd comp_0_an3v0x2_1_zn comp_0_nr2v0x2_1_a mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=82p ps=42u
M1348 comp_0_an3v0x2_1_a_24_8# comp_0_an3v0x2_1_a mux_0_gnd mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1349 comp_0_an3v0x2_1_a_31_8# comp_0_an3v0x2_2_b comp_0_an3v0x2_1_a_24_8# mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1350 comp_0_an3v0x2_1_zn mux_0_a2 comp_0_an3v0x2_1_a_31_8# mux_0_gnd nfet w=17u l=2u
+  ad=97p pd=48u as=0p ps=0u
M1351 comp_0_nr3v0x2_0_a_13_39# comp_0_an3v0x2_2_z comp_0_nr3v0x2_0_z comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=135p pd=64u as=377p ps=138u
M1352 comp_0_nr3v0x2_0_a_20_39# comp_0_an3v0x2_0_z comp_0_nr3v0x2_0_a_13_39# comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1353 mux_0_vdd comp_0_nr3v0x2_0_a comp_0_nr3v0x2_0_a_20_39# comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1354 comp_0_nr3v0x2_0_a_37_39# comp_0_nr3v0x2_0_a mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1355 comp_0_nr3v0x2_0_a_44_39# comp_0_an3v0x2_0_z comp_0_nr3v0x2_0_a_37_39# comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1356 comp_0_nr3v0x2_0_z comp_0_an3v0x2_2_z comp_0_nr3v0x2_0_a_44_39# comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1357 comp_0_nr3v0x2_0_a_61_39# comp_0_an3v0x2_2_z comp_0_nr3v0x2_0_z comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1358 comp_0_nr3v0x2_0_a_68_39# comp_0_an3v0x2_0_z comp_0_nr3v0x2_0_a_61_39# comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1359 mux_0_vdd comp_0_nr3v0x2_0_a comp_0_nr3v0x2_0_a_68_39# comp_0_an3v0x2_2_w_n4_32# pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1360 mux_0_gnd comp_0_an3v0x2_2_z comp_0_nr3v0x2_0_z mux_0_gnd nfet w=15u l=2u
+  ad=0p pd=0u as=207p ps=90u
M1361 comp_0_nr3v0x2_0_z comp_0_an3v0x2_0_z mux_0_gnd mux_0_gnd nfet w=15u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1362 mux_0_gnd comp_0_nr3v0x2_0_a comp_0_nr3v0x2_0_z mux_0_gnd nfet w=15u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1363 mux_0_vdd comp_0_an3v0x2_2_zn comp_0_an3v0x2_2_z comp_0_an3v0x2_2_w_n4_32# pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1364 comp_0_an3v0x2_2_zn mux_0_a0 mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=17u l=2u
+  ad=233p pd=98u as=0p ps=0u
M1365 mux_0_vdd comp_0_an3v0x2_2_b comp_0_an3v0x2_2_zn comp_0_an3v0x2_2_w_n4_32# pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1366 comp_0_an3v0x2_2_zn mux_0_a2 mux_0_vdd comp_0_an3v0x2_2_w_n4_32# pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1367 mux_0_gnd comp_0_an3v0x2_2_zn comp_0_an3v0x2_2_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=82p ps=42u
M1368 comp_0_an3v0x2_2_a_24_8# mux_0_a0 mux_0_gnd mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1369 comp_0_an3v0x2_2_a_31_8# comp_0_an3v0x2_2_b comp_0_an3v0x2_2_a_24_8# mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1370 comp_0_an3v0x2_2_zn mux_0_a2 comp_0_an3v0x2_2_a_31_8# mux_0_gnd nfet w=17u l=2u
+  ad=97p pd=48u as=0p ps=0u
M1371 comp_0_nr2v0x2_1_a_11_39# comp_0_nr2v0x2_1_a mux_0_vdd mux_0_vdd pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1372 comp_0_nd3v0x2_0_c comp_0_an3v0x2_3_z comp_0_nr2v0x2_1_a_11_39# mux_0_vdd pfet w=27u l=2u
+  ad=216p pd=70u as=0p ps=0u
M1373 comp_0_nr2v0x2_1_a_28_39# comp_0_an3v0x2_3_z comp_0_nd3v0x2_0_c mux_0_vdd pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1374 mux_0_vdd comp_0_nr2v0x2_1_a comp_0_nr2v0x2_1_a_28_39# mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1375 comp_0_nd3v0x2_0_c comp_0_nr2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=15u l=2u
+  ad=120p pd=46u as=0p ps=0u
M1376 mux_0_gnd comp_0_an3v0x2_3_z comp_0_nd3v0x2_0_c mux_0_gnd nfet w=15u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1377 mux_0_vdd comp_0_an3v0x2_3_zn comp_0_an3v0x2_3_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1378 comp_0_an3v0x2_3_zn comp_0_an2v0x2_0_b mux_0_vdd mux_0_vdd pfet w=17u l=2u
+  ad=233p pd=98u as=0p ps=0u
M1379 mux_0_vdd mux_0_a1 comp_0_an3v0x2_3_zn mux_0_vdd pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1380 comp_0_an3v0x2_3_zn mux_0_a0 mux_0_vdd mux_0_vdd pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1381 mux_0_gnd comp_0_an3v0x2_3_zn comp_0_an3v0x2_3_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=82p ps=42u
M1382 comp_0_an3v0x2_3_a_24_8# comp_0_an2v0x2_0_b mux_0_gnd mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1383 comp_0_an3v0x2_3_a_31_8# mux_0_a1 comp_0_an3v0x2_3_a_24_8# mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1384 comp_0_an3v0x2_3_zn mux_0_a0 comp_0_an3v0x2_3_a_31_8# mux_0_gnd nfet w=17u l=2u
+  ad=97p pd=48u as=0p ps=0u
M1385 mux_0_vdd comp_0_an3v0x2_0_zn comp_0_an3v0x2_0_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1386 comp_0_an3v0x2_0_zn comp_0_an3v0x2_1_a mux_0_vdd mux_0_vdd pfet w=17u l=2u
+  ad=233p pd=98u as=0p ps=0u
M1387 mux_0_vdd mux_0_a1 comp_0_an3v0x2_0_zn mux_0_vdd pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1388 comp_0_an3v0x2_0_zn comp_0_an2v0x2_0_b mux_0_vdd mux_0_vdd pfet w=17u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1389 mux_0_gnd comp_0_an3v0x2_0_zn comp_0_an3v0x2_0_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=82p ps=42u
M1390 comp_0_an3v0x2_0_a_24_8# comp_0_an3v0x2_1_a mux_0_gnd mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1391 comp_0_an3v0x2_0_a_31_8# mux_0_a1 comp_0_an3v0x2_0_a_24_8# mux_0_gnd nfet w=17u l=2u
+  ad=85p pd=44u as=0p ps=0u
M1392 comp_0_an3v0x2_0_zn comp_0_an2v0x2_0_b comp_0_an3v0x2_0_a_31_8# mux_0_gnd nfet w=17u l=2u
+  ad=97p pd=48u as=0p ps=0u
M1393 mux_0_vdd comp_0_an2v0x2_0_zn comp_0_nr3v0x2_0_a mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1394 comp_0_an2v0x2_0_zn mux_0_a2 mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1395 mux_0_vdd comp_0_an2v0x2_0_b comp_0_an2v0x2_0_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1396 mux_0_gnd comp_0_an2v0x2_0_zn comp_0_nr3v0x2_0_a mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1397 comp_0_an2v0x2_0_a_24_13# mux_0_a2 mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1398 comp_0_an2v0x2_0_zn comp_0_an2v0x2_0_b comp_0_an2v0x2_0_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1399 comp_0_nr2v0x2_0_a_11_39# comp_0_an2v0x2_3_z mux_0_vdd mux_0_vdd pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1400 comp_0_nd3v0x2_0_a comp_0_an2v0x2_1_z comp_0_nr2v0x2_0_a_11_39# mux_0_vdd pfet w=27u l=2u
+  ad=216p pd=70u as=0p ps=0u
M1401 comp_0_nr2v0x2_0_a_28_39# comp_0_an2v0x2_1_z comp_0_nd3v0x2_0_a mux_0_vdd pfet w=27u l=2u
+  ad=135p pd=64u as=0p ps=0u
M1402 mux_0_vdd comp_0_an2v0x2_3_z comp_0_nr2v0x2_0_a_28_39# mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1403 comp_0_nd3v0x2_0_a comp_0_an2v0x2_3_z mux_0_gnd mux_0_gnd nfet w=15u l=2u
+  ad=120p pd=46u as=0p ps=0u
M1404 mux_0_gnd comp_0_an2v0x2_1_z comp_0_nd3v0x2_0_a mux_0_gnd nfet w=15u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1405 mux_0_vdd comp_0_or3v0x2_1_zn comp_0_an2v0x2_3_b mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1406 comp_0_or3v0x2_1_a_24_38# comp_0_an3v0x2_2_b mux_0_vdd mux_0_vdd pfet w=22u l=2u
+  ad=110p pd=54u as=0p ps=0u
M1407 comp_0_or3v0x2_1_a_31_38# comp_0_an3v0x2_1_a comp_0_or3v0x2_1_a_24_38# mux_0_vdd pfet w=22u l=2u
+  ad=110p pd=54u as=0p ps=0u
M1408 comp_0_or3v0x2_1_zn mux_0_a0 comp_0_or3v0x2_1_a_31_38# mux_0_vdd pfet w=22u l=2u
+  ad=167p pd=60u as=0p ps=0u
M1409 comp_0_or3v0x2_1_a_48_38# mux_0_a0 comp_0_or3v0x2_1_zn mux_0_vdd pfet w=19u l=2u
+  ad=95p pd=48u as=0p ps=0u
M1410 comp_0_or3v0x2_1_a_55_38# comp_0_an3v0x2_1_a comp_0_or3v0x2_1_a_48_38# mux_0_vdd pfet w=19u l=2u
+  ad=95p pd=48u as=0p ps=0u
M1411 mux_0_vdd comp_0_an3v0x2_2_b comp_0_or3v0x2_1_a_55_38# mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1412 mux_0_gnd comp_0_or3v0x2_1_zn comp_0_an2v0x2_3_b mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1413 comp_0_or3v0x2_1_zn comp_0_an3v0x2_2_b mux_0_gnd mux_0_gnd nfet w=8u l=2u
+  ad=116p pd=62u as=0p ps=0u
M1414 mux_0_gnd comp_0_an3v0x2_1_a comp_0_or3v0x2_1_zn mux_0_gnd nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1415 comp_0_or3v0x2_1_zn mux_0_a0 mux_0_gnd mux_0_gnd nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1416 mux_0_vdd comp_0_an2v0x2_1_zn comp_0_an2v0x2_1_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1417 comp_0_an2v0x2_1_zn comp_0_an2v0x2_4_z mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1418 mux_0_vdd comp_0_an2v0x2_1_b comp_0_an2v0x2_1_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1419 mux_0_gnd comp_0_an2v0x2_1_zn comp_0_an2v0x2_1_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1420 comp_0_an2v0x2_1_a_24_13# comp_0_an2v0x2_4_z mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1421 comp_0_an2v0x2_1_zn comp_0_an2v0x2_1_b comp_0_an2v0x2_1_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1422 mux_0_vdd comp_0_an2v0x2_4_zn comp_0_an2v0x2_4_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1423 comp_0_an2v0x2_4_zn comp_0_an2v0x2_0_b mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1424 mux_0_vdd comp_0_an3v0x2_2_b comp_0_an2v0x2_4_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1425 mux_0_gnd comp_0_an2v0x2_4_zn comp_0_an2v0x2_4_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1426 comp_0_an2v0x2_4_a_24_13# comp_0_an2v0x2_0_b mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1427 comp_0_an2v0x2_4_zn comp_0_an3v0x2_2_b comp_0_an2v0x2_4_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1428 comp_0_an3v0x2_2_b mux_0_b1 mux_0_vdd mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1429 mux_0_vdd mux_0_b1 comp_0_an3v0x2_2_b mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1430 comp_0_an3v0x2_2_b mux_0_b1 mux_0_gnd mux_0_gnd nfet w=17u l=2u
+  ad=118p pd=50u as=0p ps=0u
M1431 mux_0_gnd mux_0_b1 comp_0_an3v0x2_2_b mux_0_gnd nfet w=11u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1432 mux_0_vdd comp_0_an2v0x2_3_zn comp_0_an2v0x2_3_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1433 comp_0_an2v0x2_3_zn comp_0_an2v0x2_2_z mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1434 mux_0_vdd comp_0_an2v0x2_3_b comp_0_an2v0x2_3_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1435 mux_0_gnd comp_0_an2v0x2_3_zn comp_0_an2v0x2_3_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1436 comp_0_an2v0x2_3_a_24_13# comp_0_an2v0x2_2_z mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1437 comp_0_an2v0x2_3_zn comp_0_an2v0x2_3_b comp_0_an2v0x2_3_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1438 mux_0_vdd comp_0_an2v0x2_2_zn comp_0_an2v0x2_2_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1439 comp_0_an2v0x2_2_zn mux_0_a2 mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1440 mux_0_vdd mux_0_a1 comp_0_an2v0x2_2_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1441 mux_0_gnd comp_0_an2v0x2_2_zn comp_0_an2v0x2_2_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1442 comp_0_an2v0x2_2_a_24_13# mux_0_a2 mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1443 comp_0_an2v0x2_2_zn mux_0_a1 comp_0_an2v0x2_2_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1444 mux_0_vdd comp_0_or3v0x2_0_zn comp_0_an2v0x2_1_b mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1445 comp_0_or3v0x2_0_a_24_38# mux_0_a1 mux_0_vdd mux_0_vdd pfet w=22u l=2u
+  ad=110p pd=54u as=0p ps=0u
M1446 comp_0_or3v0x2_0_a_31_38# mux_0_a0 comp_0_or3v0x2_0_a_24_38# mux_0_vdd pfet w=22u l=2u
+  ad=110p pd=54u as=0p ps=0u
M1447 comp_0_or3v0x2_0_zn comp_0_an3v0x2_1_a comp_0_or3v0x2_0_a_31_38# mux_0_vdd pfet w=22u l=2u
+  ad=167p pd=60u as=0p ps=0u
M1448 comp_0_or3v0x2_0_a_48_38# comp_0_an3v0x2_1_a comp_0_or3v0x2_0_zn mux_0_vdd pfet w=19u l=2u
+  ad=95p pd=48u as=0p ps=0u
M1449 comp_0_or3v0x2_0_a_55_38# mux_0_a0 comp_0_or3v0x2_0_a_48_38# mux_0_vdd pfet w=19u l=2u
+  ad=95p pd=48u as=0p ps=0u
M1450 mux_0_vdd mux_0_a1 comp_0_or3v0x2_0_a_55_38# mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1451 mux_0_gnd comp_0_or3v0x2_0_zn comp_0_an2v0x2_1_b mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1452 comp_0_or3v0x2_0_zn mux_0_a1 mux_0_gnd mux_0_gnd nfet w=8u l=2u
+  ad=116p pd=62u as=0p ps=0u
M1453 mux_0_gnd mux_0_a0 comp_0_or3v0x2_0_zn mux_0_gnd nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1454 comp_0_or3v0x2_0_zn comp_0_an3v0x2_1_a mux_0_gnd mux_0_gnd nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1455 comp_0_an3v0x2_1_a mux_0_b0 mux_0_vdd mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1456 mux_0_vdd mux_0_b0 comp_0_an3v0x2_1_a mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1457 comp_0_an3v0x2_1_a mux_0_b0 mux_0_gnd mux_0_gnd nfet w=17u l=2u
+  ad=118p pd=50u as=0p ps=0u
M1458 mux_0_gnd mux_0_b0 comp_0_an3v0x2_1_a mux_0_gnd nfet w=11u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1459 comp_0_an2v0x2_0_b mux_0_b2 mux_0_vdd mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1460 mux_0_vdd mux_0_b2 comp_0_an2v0x2_0_b mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1461 comp_0_an2v0x2_0_b mux_0_b2 mux_0_gnd mux_0_gnd nfet w=17u l=2u
+  ad=118p pd=50u as=0p ps=0u
M1462 mux_0_gnd mux_0_b2 comp_0_an2v0x2_0_b mux_0_gnd nfet w=11u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1463 mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_2_zn mux_0_b2 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1464 totdiff3_1_mux_0_mxn2v0x1_2_a_21_50# totdiff3_1_mux_0_a2 mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1465 totdiff3_1_mux_0_mxn2v0x1_2_zn totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_2_a_21_50# totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1466 totdiff3_1_mux_0_mxn2v0x1_2_a_38_50# totdiff3_1_mux_0_mxn2v0x1_2_sn totdiff3_1_mux_0_mxn2v0x1_2_zn totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1467 mux_0_vdd totdiff3_1_mux_0_b2 totdiff3_1_mux_0_mxn2v0x1_2_a_38_50# totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1468 totdiff3_1_mux_0_mxn2v0x1_2_sn totdiff3_1_mux_0_s mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1469 mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_2_zn mux_0_b2 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1470 totdiff3_1_mux_0_mxn2v0x1_2_a_21_12# totdiff3_1_mux_0_a2 mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1471 totdiff3_1_mux_0_mxn2v0x1_2_zn totdiff3_1_mux_0_mxn2v0x1_2_sn totdiff3_1_mux_0_mxn2v0x1_2_a_21_12# totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1472 totdiff3_1_mux_0_mxn2v0x1_2_a_38_12# totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_2_zn totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1473 mux_0_gnd totdiff3_1_mux_0_b2 totdiff3_1_mux_0_mxn2v0x1_2_a_38_12# totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1474 totdiff3_1_mux_0_mxn2v0x1_2_sn totdiff3_1_mux_0_s mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1475 mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_1_zn mux_0_b1 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1476 totdiff3_1_mux_0_mxn2v0x1_1_a_21_50# totdiff3_1_mux_0_a1 mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1477 totdiff3_1_mux_0_mxn2v0x1_1_zn totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_1_a_21_50# totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1478 totdiff3_1_mux_0_mxn2v0x1_1_a_38_50# totdiff3_1_mux_0_mxn2v0x1_1_sn totdiff3_1_mux_0_mxn2v0x1_1_zn totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1479 mux_0_vdd totdiff3_1_mux_0_b1 totdiff3_1_mux_0_mxn2v0x1_1_a_38_50# totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1480 totdiff3_1_mux_0_mxn2v0x1_1_sn totdiff3_1_mux_0_s mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1481 mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_1_zn mux_0_b1 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1482 totdiff3_1_mux_0_mxn2v0x1_1_a_21_12# totdiff3_1_mux_0_a1 mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1483 totdiff3_1_mux_0_mxn2v0x1_1_zn totdiff3_1_mux_0_mxn2v0x1_1_sn totdiff3_1_mux_0_mxn2v0x1_1_a_21_12# totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1484 totdiff3_1_mux_0_mxn2v0x1_1_a_38_12# totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_1_zn totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1485 mux_0_gnd totdiff3_1_mux_0_b1 totdiff3_1_mux_0_mxn2v0x1_1_a_38_12# totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1486 totdiff3_1_mux_0_mxn2v0x1_1_sn totdiff3_1_mux_0_s mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1487 mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_0_zn mux_0_b0 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1488 totdiff3_1_mux_0_mxn2v0x1_0_a_21_50# totdiff3_1_mux_0_a0 mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1489 totdiff3_1_mux_0_mxn2v0x1_0_zn totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_0_a_21_50# totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1490 totdiff3_1_mux_0_mxn2v0x1_0_a_38_50# totdiff3_1_mux_0_mxn2v0x1_0_sn totdiff3_1_mux_0_mxn2v0x1_0_zn totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1491 mux_0_vdd totdiff3_1_mux_0_b0 totdiff3_1_mux_0_mxn2v0x1_0_a_38_50# totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1492 totdiff3_1_mux_0_mxn2v0x1_0_sn totdiff3_1_mux_0_s mux_0_vdd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1493 mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_0_zn mux_0_b0 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1494 totdiff3_1_mux_0_mxn2v0x1_0_a_21_12# totdiff3_1_mux_0_a0 mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1495 totdiff3_1_mux_0_mxn2v0x1_0_zn totdiff3_1_mux_0_mxn2v0x1_0_sn totdiff3_1_mux_0_mxn2v0x1_0_a_21_12# totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1496 totdiff3_1_mux_0_mxn2v0x1_0_a_38_12# totdiff3_1_mux_0_s totdiff3_1_mux_0_mxn2v0x1_0_zn totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1497 mux_0_gnd totdiff3_1_mux_0_b0 totdiff3_1_mux_0_mxn2v0x1_0_a_38_12# totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1498 totdiff3_1_mux_0_mxn2v0x1_0_sn totdiff3_1_mux_0_s mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1499 mux_0_vdd totdiff3_1_diff2_2_an2v0x2_2_zn totdiff3_1_diff2_2_an2v0x2_2_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1500 totdiff3_1_diff2_2_an2v0x2_2_zn totdiff3_1_diff2_2_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1501 mux_0_vdd totdiff3_1_diff2_2_in_2c totdiff3_1_diff2_2_an2v0x2_2_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1502 mux_0_gnd totdiff3_1_diff2_2_an2v0x2_2_zn totdiff3_1_diff2_2_an2v0x2_2_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1503 totdiff3_1_diff2_2_an2v0x2_2_a_24_13# totdiff3_1_diff2_2_an2v0x2_2_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1504 totdiff3_1_diff2_2_an2v0x2_2_zn totdiff3_1_diff2_2_in_2c totdiff3_1_diff2_2_an2v0x2_2_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1505 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_mux_0_b2 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1506 totdiff3_1_mux_0_b2 totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_diff2_2_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1507 totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_mux_0_b2 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1508 totdiff3_1_mux_0_b2 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_diff2_2_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1509 totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_diff2_2_in_2c mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1510 mux_0_vdd totdiff3_1_diff2_2_in_2c totdiff3_1_diff2_2_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1511 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_diff2_2_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1512 mux_0_vdd totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_1_diff2_2_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1513 totdiff3_1_diff2_2_xor2v2x2_0_a_13_13# totdiff3_1_diff2_2_xor2v2x2_0_an mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1514 totdiff3_1_mux_0_b2 totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_diff2_2_xor2v2x2_0_a_13_13# mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1515 totdiff3_1_diff2_2_xor2v2x2_0_a_30_13# totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_mux_0_b2 mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1516 mux_0_gnd totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_diff2_2_xor2v2x2_0_a_30_13# mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1517 totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_diff2_2_in_2c mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1518 totdiff3_1_mux_0_b2 totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_1_diff2_2_xor2v2x2_0_bn mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1519 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_diff2_2_in_2c totdiff3_1_mux_0_b2 mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1520 mux_0_gnd totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_1_diff2_2_xor2v2x2_0_an mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1521 totdiff3_1_mux_0_s totdiff3_1_diff2_2_or2v0x3_0_zn mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1522 mux_0_vdd totdiff3_1_diff2_2_or2v0x3_0_zn totdiff3_1_mux_0_s mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1523 totdiff3_1_diff2_2_or2v0x3_0_a_31_39# totdiff3_1_diff2_2_an2v0x2_1_z mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1524 totdiff3_1_diff2_2_or2v0x3_0_zn totdiff3_1_diff2_2_an2v0x2_0_z totdiff3_1_diff2_2_or2v0x3_0_a_31_39# mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1525 totdiff3_1_diff2_2_or2v0x3_0_a_48_39# totdiff3_1_diff2_2_an2v0x2_0_z totdiff3_1_diff2_2_or2v0x3_0_zn mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1526 mux_0_vdd totdiff3_1_diff2_2_an2v0x2_1_z totdiff3_1_diff2_2_or2v0x3_0_a_48_39# mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1527 mux_0_gnd totdiff3_1_diff2_2_or2v0x3_0_zn totdiff3_1_mux_0_s mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1528 totdiff3_1_diff2_2_or2v0x3_0_zn totdiff3_1_diff2_2_an2v0x2_1_z mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1529 mux_0_gnd totdiff3_1_diff2_2_an2v0x2_0_z totdiff3_1_diff2_2_or2v0x3_0_zn mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1530 mux_0_vdd totdiff3_1_diff2_2_an2v0x2_1_zn totdiff3_1_diff2_2_an2v0x2_1_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1531 totdiff3_1_diff2_2_an2v0x2_1_zn totdiff3_1_diff2_2_an2v0x2_1_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1532 mux_0_vdd totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_an2v0x2_1_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1533 mux_0_gnd totdiff3_1_diff2_2_an2v0x2_1_zn totdiff3_1_diff2_2_an2v0x2_1_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1534 totdiff3_1_diff2_2_an2v0x2_1_a_24_13# totdiff3_1_diff2_2_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1535 totdiff3_1_diff2_2_an2v0x2_1_zn totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_an2v0x2_1_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1536 mux_0_vdd totdiff3_1_diff2_2_an2v0x2_0_zn totdiff3_1_diff2_2_an2v0x2_0_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1537 totdiff3_1_diff2_2_an2v0x2_0_zn totdiff3_1_diff2_2_in_c mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1538 mux_0_vdd totdiff3_1_diff2_2_an2v0x2_0_b totdiff3_1_diff2_2_an2v0x2_0_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1539 mux_0_gnd totdiff3_1_diff2_2_an2v0x2_0_zn totdiff3_1_diff2_2_an2v0x2_0_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1540 totdiff3_1_diff2_2_an2v0x2_0_a_24_13# totdiff3_1_diff2_2_in_c mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1541 totdiff3_1_diff2_2_an2v0x2_0_zn totdiff3_1_diff2_2_an2v0x2_0_b totdiff3_1_diff2_2_an2v0x2_0_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1542 mux_0_vdd totdiff3_1_diff2_2_xnr2v8x05_0_zn totdiff3_1_diff2_2_an2v0x2_0_b mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1543 totdiff3_1_diff2_2_xnr2v8x05_0_an totdiff3_1_diff2_2_in_a mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1544 totdiff3_1_diff2_2_xnr2v8x05_0_zn totdiff3_1_diff2_2_xnr2v8x05_0_bn totdiff3_1_diff2_2_xnr2v8x05_0_an mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1545 totdiff3_1_diff2_2_xnr2v8x05_0_ai totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_xnr2v8x05_0_zn mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1546 mux_0_vdd totdiff3_1_diff2_2_xnr2v8x05_0_an totdiff3_1_diff2_2_xnr2v8x05_0_ai mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1547 totdiff3_1_diff2_2_xnr2v8x05_0_bn totdiff3_1_diff2_2_in_b mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1548 mux_0_gnd totdiff3_1_diff2_2_xnr2v8x05_0_zn totdiff3_1_diff2_2_an2v0x2_0_b mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1549 totdiff3_1_diff2_2_xnr2v8x05_0_an totdiff3_1_diff2_2_in_a mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1550 totdiff3_1_diff2_2_xnr2v8x05_0_zn totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_xnr2v8x05_0_an mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1551 totdiff3_1_diff2_2_xnr2v8x05_0_ai totdiff3_1_diff2_2_xnr2v8x05_0_bn totdiff3_1_diff2_2_xnr2v8x05_0_zn mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1552 mux_0_gnd totdiff3_1_diff2_2_xnr2v8x05_0_an totdiff3_1_diff2_2_xnr2v8x05_0_ai mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1553 totdiff3_1_diff2_2_xnr2v8x05_0_bn totdiff3_1_diff2_2_in_b mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1554 totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_1_mux_0_a2 mux_0_vdd mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1555 mux_0_vdd totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_an2v0x2_2_a mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1556 totdiff3_1_diff2_2_an2v0x2_2_a totdiff3_1_mux_0_a2 mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1557 mux_0_gnd totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_an2v0x2_2_a mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1558 totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_mux_0_a2 mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1559 totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_xor3v1x2_0_cn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1560 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_mux_0_a2 mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1561 totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_diff2_2_xor3v1x2_0_zn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1562 totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_diff2_2_in_c mux_0_vdd mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1563 mux_0_vdd totdiff3_1_diff2_2_in_c totdiff3_1_diff2_2_xor3v1x2_0_cn mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1564 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_xor3v1x2_0_iz mux_0_vdd mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1565 mux_0_vdd totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_1_diff2_2_xor3v1x2_0_zn mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1566 totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_1_diff2_2_xor3v1x2_0_bn mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1567 totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_1_diff2_2_xor3v1x2_0_bn totdiff3_1_diff2_2_xor3v1x2_0_iz mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1568 mux_0_vdd totdiff3_1_diff2_2_in_a totdiff3_1_diff2_2_an2v0x2_1_a mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1569 totdiff3_1_diff2_2_xor3v1x2_0_bn totdiff3_1_diff2_2_in_b mux_0_vdd mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1570 mux_0_vdd totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_xor3v1x2_0_bn mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1571 totdiff3_1_diff2_2_xor3v1x2_0_a_11_12# totdiff3_1_diff2_2_xor3v1x2_0_cn mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1572 totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_xor3v1x2_0_a_11_12# mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1573 totdiff3_1_diff2_2_xor3v1x2_0_a_28_12# totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_mux_0_a2 mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1574 mux_0_gnd totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_diff2_2_xor3v1x2_0_a_28_12# mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1575 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_xor3v1x2_0_iz mux_0_gnd mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1576 totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_in_c totdiff3_1_diff2_2_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1577 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_in_c totdiff3_1_mux_0_a2 mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1578 mux_0_gnd totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_1_diff2_2_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1579 totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_diff2_2_in_c mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1580 mux_0_gnd totdiff3_1_diff2_2_in_c totdiff3_1_diff2_2_xor3v1x2_0_cn mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1581 totdiff3_1_diff2_2_xor3v1x2_0_a_115_7# totdiff3_1_diff2_2_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1582 totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_1_diff2_2_xor3v1x2_0_bn totdiff3_1_diff2_2_xor3v1x2_0_a_115_7# mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1583 totdiff3_1_diff2_2_an2v0x2_1_a totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_xor3v1x2_0_iz mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1584 mux_0_gnd totdiff3_1_diff2_2_in_a totdiff3_1_diff2_2_an2v0x2_1_a mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1585 totdiff3_1_diff2_2_xor3v1x2_0_bn totdiff3_1_diff2_2_in_b mux_0_gnd mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1586 mux_0_vdd totdiff3_1_diff2_1_an2v0x2_2_zn totdiff3_1_diff2_2_in_2c mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1587 totdiff3_1_diff2_1_an2v0x2_2_zn totdiff3_1_diff2_1_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1588 mux_0_vdd totdiff3_1_diff2_1_in_2c totdiff3_1_diff2_1_an2v0x2_2_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1589 mux_0_gnd totdiff3_1_diff2_1_an2v0x2_2_zn totdiff3_1_diff2_2_in_2c mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1590 totdiff3_1_diff2_1_an2v0x2_2_a_24_13# totdiff3_1_diff2_1_an2v0x2_2_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1591 totdiff3_1_diff2_1_an2v0x2_2_zn totdiff3_1_diff2_1_in_2c totdiff3_1_diff2_1_an2v0x2_2_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1592 totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_mux_0_b1 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1593 totdiff3_1_mux_0_b1 totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_diff2_1_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1594 totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_1_mux_0_b1 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1595 totdiff3_1_mux_0_b1 totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_1_diff2_1_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1596 totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_diff2_1_in_2c mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1597 mux_0_vdd totdiff3_1_diff2_1_in_2c totdiff3_1_diff2_1_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1598 totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_1_diff2_1_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1599 mux_0_vdd totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_1_diff2_1_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1600 totdiff3_1_diff2_1_xor2v2x2_0_a_13_13# totdiff3_1_diff2_1_xor2v2x2_0_an mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1601 totdiff3_1_mux_0_b1 totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_diff2_1_xor2v2x2_0_a_13_13# mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1602 totdiff3_1_diff2_1_xor2v2x2_0_a_30_13# totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_mux_0_b1 mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1603 mux_0_gnd totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_1_diff2_1_xor2v2x2_0_a_30_13# mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1604 totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_diff2_1_in_2c mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1605 totdiff3_1_mux_0_b1 totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_1_diff2_1_xor2v2x2_0_bn mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1606 totdiff3_1_diff2_1_xor2v2x2_0_an totdiff3_1_diff2_1_in_2c totdiff3_1_mux_0_b1 mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1607 mux_0_gnd totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_1_diff2_1_xor2v2x2_0_an mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1608 totdiff3_1_diff2_2_in_c totdiff3_1_diff2_1_or2v0x3_0_zn mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1609 mux_0_vdd totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_1_diff2_2_in_c mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1610 totdiff3_1_diff2_1_or2v0x3_0_a_31_39# totdiff3_1_diff2_1_an2v0x2_1_z mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1611 totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_1_diff2_1_an2v0x2_0_z totdiff3_1_diff2_1_or2v0x3_0_a_31_39# mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1612 totdiff3_1_diff2_1_or2v0x3_0_a_48_39# totdiff3_1_diff2_1_an2v0x2_0_z totdiff3_1_diff2_1_or2v0x3_0_zn mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1613 mux_0_vdd totdiff3_1_diff2_1_an2v0x2_1_z totdiff3_1_diff2_1_or2v0x3_0_a_48_39# mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1614 mux_0_gnd totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_1_diff2_2_in_c mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1615 totdiff3_1_diff2_1_or2v0x3_0_zn totdiff3_1_diff2_1_an2v0x2_1_z mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1616 mux_0_gnd totdiff3_1_diff2_1_an2v0x2_0_z totdiff3_1_diff2_1_or2v0x3_0_zn mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1617 mux_0_vdd totdiff3_1_diff2_1_an2v0x2_1_zn totdiff3_1_diff2_1_an2v0x2_1_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1618 totdiff3_1_diff2_1_an2v0x2_1_zn totdiff3_1_diff2_1_an2v0x2_1_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1619 mux_0_vdd totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_an2v0x2_1_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1620 mux_0_gnd totdiff3_1_diff2_1_an2v0x2_1_zn totdiff3_1_diff2_1_an2v0x2_1_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1621 totdiff3_1_diff2_1_an2v0x2_1_a_24_13# totdiff3_1_diff2_1_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1622 totdiff3_1_diff2_1_an2v0x2_1_zn totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_an2v0x2_1_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1623 mux_0_vdd totdiff3_1_diff2_1_an2v0x2_0_zn totdiff3_1_diff2_1_an2v0x2_0_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1624 totdiff3_1_diff2_1_an2v0x2_0_zn totdiff3_1_diff2_1_in_c mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1625 mux_0_vdd totdiff3_1_diff2_1_an2v0x2_0_b totdiff3_1_diff2_1_an2v0x2_0_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1626 mux_0_gnd totdiff3_1_diff2_1_an2v0x2_0_zn totdiff3_1_diff2_1_an2v0x2_0_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1627 totdiff3_1_diff2_1_an2v0x2_0_a_24_13# totdiff3_1_diff2_1_in_c mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1628 totdiff3_1_diff2_1_an2v0x2_0_zn totdiff3_1_diff2_1_an2v0x2_0_b totdiff3_1_diff2_1_an2v0x2_0_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1629 mux_0_vdd totdiff3_1_diff2_1_xnr2v8x05_0_zn totdiff3_1_diff2_1_an2v0x2_0_b mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1630 totdiff3_1_diff2_1_xnr2v8x05_0_an totdiff3_1_diff2_1_in_a mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1631 totdiff3_1_diff2_1_xnr2v8x05_0_zn totdiff3_1_diff2_1_xnr2v8x05_0_bn totdiff3_1_diff2_1_xnr2v8x05_0_an mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1632 totdiff3_1_diff2_1_xnr2v8x05_0_ai totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_xnr2v8x05_0_zn mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1633 mux_0_vdd totdiff3_1_diff2_1_xnr2v8x05_0_an totdiff3_1_diff2_1_xnr2v8x05_0_ai mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1634 totdiff3_1_diff2_1_xnr2v8x05_0_bn totdiff3_1_diff2_1_in_b mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1635 mux_0_gnd totdiff3_1_diff2_1_xnr2v8x05_0_zn totdiff3_1_diff2_1_an2v0x2_0_b mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1636 totdiff3_1_diff2_1_xnr2v8x05_0_an totdiff3_1_diff2_1_in_a mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1637 totdiff3_1_diff2_1_xnr2v8x05_0_zn totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_xnr2v8x05_0_an mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1638 totdiff3_1_diff2_1_xnr2v8x05_0_ai totdiff3_1_diff2_1_xnr2v8x05_0_bn totdiff3_1_diff2_1_xnr2v8x05_0_zn mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1639 mux_0_gnd totdiff3_1_diff2_1_xnr2v8x05_0_an totdiff3_1_diff2_1_xnr2v8x05_0_ai mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1640 totdiff3_1_diff2_1_xnr2v8x05_0_bn totdiff3_1_diff2_1_in_b mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1641 totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_1_mux_0_a1 mux_0_vdd mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1642 mux_0_vdd totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_an2v0x2_2_a mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1643 totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_1_mux_0_a1 mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1644 mux_0_gnd totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_an2v0x2_2_a mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1645 totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_mux_0_a1 mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1646 totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_xor3v1x2_0_cn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1647 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_mux_0_a1 mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1648 totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_diff2_1_xor3v1x2_0_zn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1649 totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_diff2_1_in_c mux_0_vdd mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1650 mux_0_vdd totdiff3_1_diff2_1_in_c totdiff3_1_diff2_1_xor3v1x2_0_cn mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1651 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_xor3v1x2_0_iz mux_0_vdd mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1652 mux_0_vdd totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_1_diff2_1_xor3v1x2_0_zn mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1653 totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_1_diff2_1_xor3v1x2_0_bn mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1654 totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_1_diff2_1_xor3v1x2_0_iz mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1655 mux_0_vdd totdiff3_1_diff2_1_in_a totdiff3_1_diff2_1_an2v0x2_1_a mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1656 totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_1_diff2_1_in_b mux_0_vdd mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1657 mux_0_vdd totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_xor3v1x2_0_bn mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1658 totdiff3_1_diff2_1_xor3v1x2_0_a_11_12# totdiff3_1_diff2_1_xor3v1x2_0_cn mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1659 totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_xor3v1x2_0_a_11_12# mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1660 totdiff3_1_diff2_1_xor3v1x2_0_a_28_12# totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_mux_0_a1 mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1661 mux_0_gnd totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_diff2_1_xor3v1x2_0_a_28_12# mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1662 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_xor3v1x2_0_iz mux_0_gnd mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1663 totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_in_c totdiff3_1_diff2_1_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1664 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_in_c totdiff3_1_mux_0_a1 mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1665 mux_0_gnd totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_1_diff2_1_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1666 totdiff3_1_diff2_1_xor3v1x2_0_cn totdiff3_1_diff2_1_in_c mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1667 mux_0_gnd totdiff3_1_diff2_1_in_c totdiff3_1_diff2_1_xor3v1x2_0_cn mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1668 totdiff3_1_diff2_1_xor3v1x2_0_a_115_7# totdiff3_1_diff2_1_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1669 totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_1_diff2_1_xor3v1x2_0_a_115_7# mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1670 totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_1_diff2_1_in_b totdiff3_1_diff2_1_xor3v1x2_0_iz mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1671 mux_0_gnd totdiff3_1_diff2_1_in_a totdiff3_1_diff2_1_an2v0x2_1_a mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1672 totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_1_diff2_1_in_b mux_0_gnd mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1673 mux_0_vdd totdiff3_1_diff2_0_an2v0x2_2_zn totdiff3_1_diff2_1_in_2c mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1674 totdiff3_1_diff2_0_an2v0x2_2_zn totdiff3_1_diff2_0_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1675 mux_0_vdd mux_0_vdd totdiff3_1_diff2_0_an2v0x2_2_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1676 mux_0_gnd totdiff3_1_diff2_0_an2v0x2_2_zn totdiff3_1_diff2_1_in_2c mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1677 totdiff3_1_diff2_0_an2v0x2_2_a_24_13# totdiff3_1_diff2_0_an2v0x2_2_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1678 totdiff3_1_diff2_0_an2v0x2_2_zn mux_0_vdd totdiff3_1_diff2_0_an2v0x2_2_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1679 totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_1_mux_0_b0 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1680 totdiff3_1_mux_0_b0 totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_1_diff2_0_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1681 totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_1_mux_0_b0 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1682 totdiff3_1_mux_0_b0 totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_1_diff2_0_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1683 totdiff3_1_diff2_0_xor2v2x2_0_bn mux_0_vdd mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1684 mux_0_vdd mux_0_vdd totdiff3_1_diff2_0_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1685 totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_1_diff2_0_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1686 mux_0_vdd totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_1_diff2_0_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1687 totdiff3_1_diff2_0_xor2v2x2_0_a_13_13# totdiff3_1_diff2_0_xor2v2x2_0_an mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1688 totdiff3_1_mux_0_b0 totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_1_diff2_0_xor2v2x2_0_a_13_13# mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1689 totdiff3_1_diff2_0_xor2v2x2_0_a_30_13# totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_1_mux_0_b0 mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1690 mux_0_gnd totdiff3_1_diff2_0_xor2v2x2_0_an totdiff3_1_diff2_0_xor2v2x2_0_a_30_13# mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1691 totdiff3_1_diff2_0_xor2v2x2_0_bn mux_0_vdd mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1692 totdiff3_1_mux_0_b0 totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_1_diff2_0_xor2v2x2_0_bn mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1693 totdiff3_1_diff2_0_xor2v2x2_0_an mux_0_vdd totdiff3_1_mux_0_b0 mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1694 mux_0_gnd totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_1_diff2_0_xor2v2x2_0_an mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1695 totdiff3_1_diff2_1_in_c totdiff3_1_diff2_0_or2v0x3_0_zn mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1696 mux_0_vdd totdiff3_1_diff2_0_or2v0x3_0_zn totdiff3_1_diff2_1_in_c mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1697 totdiff3_1_diff2_0_or2v0x3_0_a_31_39# totdiff3_1_diff2_0_an2v0x2_1_z mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1698 totdiff3_1_diff2_0_or2v0x3_0_zn totdiff3_1_diff2_0_an2v0x2_0_z totdiff3_1_diff2_0_or2v0x3_0_a_31_39# mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1699 totdiff3_1_diff2_0_or2v0x3_0_a_48_39# totdiff3_1_diff2_0_an2v0x2_0_z totdiff3_1_diff2_0_or2v0x3_0_zn mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1700 mux_0_vdd totdiff3_1_diff2_0_an2v0x2_1_z totdiff3_1_diff2_0_or2v0x3_0_a_48_39# mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1701 mux_0_gnd totdiff3_1_diff2_0_or2v0x3_0_zn totdiff3_1_diff2_1_in_c mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1702 totdiff3_1_diff2_0_or2v0x3_0_zn totdiff3_1_diff2_0_an2v0x2_1_z mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1703 mux_0_gnd totdiff3_1_diff2_0_an2v0x2_0_z totdiff3_1_diff2_0_or2v0x3_0_zn mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1704 mux_0_vdd totdiff3_1_diff2_0_an2v0x2_1_zn totdiff3_1_diff2_0_an2v0x2_1_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1705 totdiff3_1_diff2_0_an2v0x2_1_zn totdiff3_1_diff2_0_an2v0x2_1_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1706 mux_0_vdd totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_an2v0x2_1_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1707 mux_0_gnd totdiff3_1_diff2_0_an2v0x2_1_zn totdiff3_1_diff2_0_an2v0x2_1_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1708 totdiff3_1_diff2_0_an2v0x2_1_a_24_13# totdiff3_1_diff2_0_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1709 totdiff3_1_diff2_0_an2v0x2_1_zn totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_an2v0x2_1_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1710 mux_0_vdd totdiff3_1_diff2_0_an2v0x2_0_zn totdiff3_1_diff2_0_an2v0x2_0_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1711 totdiff3_1_diff2_0_an2v0x2_0_zn mux_0_gnd mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1712 mux_0_vdd totdiff3_1_diff2_0_an2v0x2_0_b totdiff3_1_diff2_0_an2v0x2_0_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1713 mux_0_gnd totdiff3_1_diff2_0_an2v0x2_0_zn totdiff3_1_diff2_0_an2v0x2_0_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1714 totdiff3_1_diff2_0_an2v0x2_0_a_24_13# mux_0_gnd mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1715 totdiff3_1_diff2_0_an2v0x2_0_zn totdiff3_1_diff2_0_an2v0x2_0_b totdiff3_1_diff2_0_an2v0x2_0_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1716 mux_0_vdd totdiff3_1_diff2_0_xnr2v8x05_0_zn totdiff3_1_diff2_0_an2v0x2_0_b mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1717 totdiff3_1_diff2_0_xnr2v8x05_0_an totdiff3_1_diff2_0_in_a mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1718 totdiff3_1_diff2_0_xnr2v8x05_0_zn totdiff3_1_diff2_0_xnr2v8x05_0_bn totdiff3_1_diff2_0_xnr2v8x05_0_an mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1719 totdiff3_1_diff2_0_xnr2v8x05_0_ai totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_xnr2v8x05_0_zn mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1720 mux_0_vdd totdiff3_1_diff2_0_xnr2v8x05_0_an totdiff3_1_diff2_0_xnr2v8x05_0_ai mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1721 totdiff3_1_diff2_0_xnr2v8x05_0_bn totdiff3_1_diff2_0_in_b mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1722 mux_0_gnd totdiff3_1_diff2_0_xnr2v8x05_0_zn totdiff3_1_diff2_0_an2v0x2_0_b mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1723 totdiff3_1_diff2_0_xnr2v8x05_0_an totdiff3_1_diff2_0_in_a mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1724 totdiff3_1_diff2_0_xnr2v8x05_0_zn totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_xnr2v8x05_0_an mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1725 totdiff3_1_diff2_0_xnr2v8x05_0_ai totdiff3_1_diff2_0_xnr2v8x05_0_bn totdiff3_1_diff2_0_xnr2v8x05_0_zn mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1726 mux_0_gnd totdiff3_1_diff2_0_xnr2v8x05_0_an totdiff3_1_diff2_0_xnr2v8x05_0_ai mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1727 totdiff3_1_diff2_0_xnr2v8x05_0_bn totdiff3_1_diff2_0_in_b mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1728 totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_1_mux_0_a0 mux_0_vdd mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1729 mux_0_vdd totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_an2v0x2_2_a mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1730 totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_1_mux_0_a0 mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1731 mux_0_gnd totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_an2v0x2_2_a mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1732 totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_mux_0_a0 mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1733 totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_diff2_0_xor3v1x2_0_cn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1734 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_1_mux_0_a0 mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1735 totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_1_diff2_0_xor3v1x2_0_zn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1736 totdiff3_1_diff2_0_xor3v1x2_0_cn mux_0_gnd mux_0_vdd mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1737 mux_0_vdd mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_cn mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1738 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_diff2_0_xor3v1x2_0_iz mux_0_vdd mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1739 mux_0_vdd totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_1_diff2_0_xor3v1x2_0_zn mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1740 totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_1_diff2_0_an2v0x2_1_a totdiff3_1_diff2_0_xor3v1x2_0_bn mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1741 totdiff3_1_diff2_0_an2v0x2_1_a totdiff3_1_diff2_0_xor3v1x2_0_bn totdiff3_1_diff2_0_xor3v1x2_0_iz mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1742 mux_0_vdd totdiff3_1_diff2_0_in_a totdiff3_1_diff2_0_an2v0x2_1_a mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1743 totdiff3_1_diff2_0_xor3v1x2_0_bn totdiff3_1_diff2_0_in_b mux_0_vdd mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1744 mux_0_vdd totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_xor3v1x2_0_bn mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1745 totdiff3_1_diff2_0_xor3v1x2_0_a_11_12# totdiff3_1_diff2_0_xor3v1x2_0_cn mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1746 totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_diff2_0_xor3v1x2_0_a_11_12# mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1747 totdiff3_1_diff2_0_xor3v1x2_0_a_28_12# totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_mux_0_a0 mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1748 mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_cn totdiff3_1_diff2_0_xor3v1x2_0_a_28_12# mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1749 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_diff2_0_xor3v1x2_0_iz mux_0_gnd mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1750 totdiff3_1_mux_0_a0 mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1751 totdiff3_1_diff2_0_xor3v1x2_0_zn mux_0_gnd totdiff3_1_mux_0_a0 mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1752 mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_1_diff2_0_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1753 totdiff3_1_diff2_0_xor3v1x2_0_cn mux_0_gnd mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1754 mux_0_gnd mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_cn mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1755 totdiff3_1_diff2_0_xor3v1x2_0_a_115_7# totdiff3_1_diff2_0_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1756 totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_1_diff2_0_xor3v1x2_0_bn totdiff3_1_diff2_0_xor3v1x2_0_a_115_7# mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1757 totdiff3_1_diff2_0_an2v0x2_1_a totdiff3_1_diff2_0_in_b totdiff3_1_diff2_0_xor3v1x2_0_iz mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1758 mux_0_gnd totdiff3_1_diff2_0_in_a totdiff3_1_diff2_0_an2v0x2_1_a mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1759 totdiff3_1_diff2_0_xor3v1x2_0_bn totdiff3_1_diff2_0_in_b mux_0_gnd mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
C0 mux_0_mxn2v0x1_0_zn mux_0_mxn2v0x1_0_w_n4_32# 9.3fF
C1 totdiff3_0_diff2_1_in_a mux_0_gnd 27.8fF
C2 totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_diff2_0_xor3v1x2_0_iz 2.4fF
C3 totdiff3_1_diff2_0_or2v0x3_0_zn mux_0_vdd 12.7fF
C4 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_1_mux_0_s 15.2fF
C5 totdiff3_0_diff2_1_an2v0x2_2_zn mux_0_vdd 8.8fF
C6 totdiff3_0_mux_0_a0 mux_0_gnd 14.9fF
C7 totdiff3_1_mux_0_mxn2v0x1_0_sn mux_0_b0 4.3fF
C8 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_mxn2v0x1_1_sn 9.3fF
C9 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_xor3v1x2_0_cn 4.5fF
C10 totdiff3_0_diff2_1_xnr2v8x05_0_zn mux_0_gnd 11.9fF
C11 totdiff3_1_mux_0_mxn2v0x1_1_zn totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 9.3fF
C12 totdiff3_0_diff2_1_an2v0x2_1_z mux_0_gnd 10.2fF
C13 totdiff3_0_diff2_1_xor2v2x2_0_an mux_0_gnd 21.6fF
C14 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# mux_0_a1 5.0fF
C15 totdiff3_1_mux_0_b0 mux_0_vdd 30.6fF
C16 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_1_mux_0_s 36.4fF
C17 totdiff3_1_diff2_1_or2v0x3_0_zn mux_0_gnd 9.0fF
C18 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_0_mux_0_s 18.7fF
C19 mux_0_b2 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# 2.3fF
C20 totdiff3_0_mux_0_b2 totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# 8.7fF
C21 mux_0_a1 mux_0_mxn2v0x1_0_w_n4_n4# 4.8fF
C22 totdiff3_0_mux_0_b0 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 8.7fF
C23 totdiff3_0_diff2_1_in_c mux_0_vdd 39.6fF
C24 totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_xor3v1x2_0_zn 4.6fF
C25 mux_0_a0 mux_0_b1 3.3fF
C26 mux_0_b2 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 6.3fF
C27 mux_0_mxn2v0x1_0_w_n4_32# mux_0_b0 6.6fF
C28 totdiff3_0_diff2_0_xnr2v8x05_0_an mux_0_gnd 6.8fF
C29 totdiff3_1_mux_0_mxn2v0x1_1_zn totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# 8.9fF
C30 comp_0_an3v0x2_2_zn mux_0_gnd 8.8fF
C31 totdiff3_0_diff2_0_xor3v1x2_0_bn mux_0_vdd 15.4fF
C32 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_1_mux_0_s 30.3fF
C33 totdiff3_0_diff2_2_xnr2v8x05_0_an mux_0_vdd 9.9fF
C34 mux_0_a1 mux_0_vdd 52.8fF
C35 totdiff3_1_diff2_0_an2v0x2_1_a mux_0_vdd 12.4fF
C36 comp_0_an2v0x2_0_zn mux_0_vdd 8.8fF
C37 totdiff3_0_diff2_2_xor3v1x2_0_bn mux_0_gnd 9.1fF
C38 totdiff3_0_diff2_2_an2v0x2_2_zn mux_0_gnd 8.9fF
C39 totdiff3_1_diff2_2_xor3v1x2_0_zn mux_0_gnd 11.9fF
C40 comp_0_an2v0x2_3_b mux_0_vdd 13.7fF
C41 comp_0_an3v0x2_1_a comp_0_an2v0x2_0_b 2.5fF
C42 totdiff3_1_diff2_2_xor2v2x2_0_bn mux_0_vdd 17.7fF
C43 comp_0_nd3v0x2_0_c mux_0_vdd 5.0fF
C44 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_1_mux_0_mxn2v0x1_0_zn 9.3fF
C45 mux_0_gnd totdiff3_1_diff2_1_xnr2v8x05_0_bn 6.7fF
C46 totdiff3_0_diff2_2_xor3v1x2_0_iz mux_0_vdd 15.8fF
C47 totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_an2v0x2_1_a 2.0fF
C48 comp_0_an3v0x2_3_z mux_0_vdd 15.4fF
C49 comp_0_an3v0x2_2_z mux_0_vdd 3.3fF
C50 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_diff2_0_xor3v1x2_0_cn 4.5fF
C51 mux_0_vdd totdiff3_1_diff2_0_xnr2v8x05_0_bn 14.4fF
C52 totdiff3_1_diff2_1_xnr2v8x05_0_an mux_0_vdd 9.9fF
C53 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_b1 10.2fF
C54 comp_0_an2v0x2_1_zn mux_0_vdd 8.8fF
C55 totdiff3_0_diff2_2_an2v0x2_0_z mux_0_gnd 12.8fF
C56 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_mxn2v0x1_2_sn 9.3fF
C57 comp_0_an3v0x2_2_w_n4_32# comp_0_nd3v0x2_0_c 5.7fF
C58 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# mux_0_gnd 78.2fF
C59 totdiff3_0_diff2_0_in_b mux_0_gnd 60.8fF
C60 totdiff3_0_diff2_0_an2v0x2_2_zn mux_0_vdd 10.3fF
C61 mux_0_vdd totdiff3_1_mux_0_b2 3.1fF
C62 totdiff3_1_diff2_1_xor3v1x2_0_iz totdiff3_1_diff2_1_xor3v1x2_0_bn 2.4fF
C63 comp_0_an3v0x2_2_w_n4_32# comp_0_an3v0x2_2_z 21.1fF
C64 totdiff3_0_diff2_2_in_a mux_0_vdd 24.6fF
C65 totdiff3_0_mux_0_s mux_0_gnd 8.3fF
C66 mux_0_b1 mux_0_vdd 14.0fF
C67 mux_0_vdd totdiff3_1_diff2_1_xor3v1x2_0_iz 15.8fF
C68 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_0_mux_0_mxn2v0x1_0_zn 9.3fF
C69 comp_0_an3v0x2_1_a mux_0_gnd 57.3fF
C70 totdiff3_0_diff2_0_in_b totdiff3_0_diff2_0_xor3v1x2_0_zn 4.3fF
C71 mux_0_gnd totdiff3_1_diff2_0_an2v0x2_2_a 25.9fF
C72 totdiff3_1_diff2_0_an2v0x2_1_z mux_0_vdd 17.9fF
C73 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_mxn2v0x1_1_zn 9.3fF
C74 totdiff3_1_diff2_1_an2v0x2_0_zn mux_0_gnd 8.9fF
C75 totdiff3_1_diff2_2_an2v0x2_0_zn mux_0_vdd 8.8fF
C76 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# mux_0_b0 2.3fF
C77 mux_0_vdd totdiff3_1_diff2_0_an2v0x2_0_z 24.6fF
C78 totdiff3_0_mux_0_b0 totdiff3_0_mux_0_mxn2v0x1_0_zn 2.7fF
C79 mux_0_s mux_0_mxn2v0x1_0_w_n4_n4# 30.3fF
C80 mux_0_mxn2v0x1_2_w_n4_n4# mux_0_b2 8.7fF
C81 mux_0_mxn2v0x1_1_w_n4_32# mux_0_b2 6.6fF
C82 totdiff3_1_diff2_2_xnr2v8x05_0_an mux_0_vdd 9.9fF
C83 mux_0_vdd totdiff3_1_diff2_0_xor3v1x2_0_zn 18.9fF
C84 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_1_mux_0_b0 8.7fF
C85 totdiff3_1_diff2_2_in_2c mux_0_vdd 33.2fF
C86 totdiff3_0_diff2_0_an2v0x2_0_zn mux_0_gnd 10.8fF
C87 mux_0_s mux_0_vdd 4.5fF
C88 mux_0_gnd totdiff3_1_diff2_2_an2v0x2_0_z 12.8fF
C89 mux_0_vdd totdiff3_1_diff2_0_xnr2v8x05_0_an 9.9fF
C90 mux_0_a1 mux_0_a2 10.0fF
C91 totdiff3_0_diff2_2_in_2c mux_0_gnd 17.8fF
C92 totdiff3_1_diff2_1_an2v0x2_1_a mux_0_vdd 12.4fF
C93 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_1_mux_0_a0 11.6fF
C94 comp_0_an3v0x2_1_a comp_0_an3v0x2_2_b 5.2fF
C95 mux_0_gnd totdiff3_1_diff2_2_an2v0x2_1_z 10.2fF
C96 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_1_mux_0_b2 8.7fF
C97 totdiff3_0_diff2_1_xor3v1x2_0_cn mux_0_gnd 18.8fF
C98 totdiff3_1_diff2_2_in_b totdiff3_1_diff2_2_xor3v1x2_0_bn 2.6fF
C99 totdiff3_0_diff2_1_an2v0x2_0_zn mux_0_gnd 8.9fF
C100 totdiff3_0_mux_0_mxn2v0x1_0_sn mux_0_a0 4.3fF
C101 totdiff3_0_mux_0_b2 totdiff3_0_mux_0_mxn2v0x1_2_zn 2.7fF
C102 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_diff2_2_in_b 4.3fF
C103 mux_0_gnd totdiff3_1_mux_0_s 8.3fF
C104 mux_0_gnd comp_0_or3v0x2_0_zn 10.9fF
C105 totdiff3_1_mux_0_b1 totdiff3_1_mux_0_a1 39.4fF
C106 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_1_mux_0_b2 6.6fF
C107 mux_0_vdd totdiff3_1_diff2_0_xor2v2x2_0_an 27.4fF
C108 comp_0_an2v0x2_3_z mux_0_vdd 9.1fF
C109 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_a2 11.6fF
C110 mux_0_s mux_0_mxn2v0x1_0_w_n4_32# 18.7fF
C111 totdiff3_1_diff2_2_an2v0x2_1_a mux_0_vdd 12.4fF
C112 comp_0_an3v0x2_2_zn comp_0_nr3v0x2_0_a 2.1fF
C113 totdiff3_0_diff2_0_an2v0x2_0_zn totdiff3_0_diff2_0_in_a 2.2fF
C114 totdiff3_1_diff2_2_in_b mux_0_vdd 50.3fF
C115 totdiff3_0_mux_0_a1 mux_0_gnd 15.3fF
C116 mux_0_b2 mux_0_gnd 11.2fF
C117 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# mux_0_b1 5.0fF
C118 mux_0_mxn2v0x1_2_w_n4_n4# mux_0_mxn2v0x1_2_zn 8.9fF
C119 mux_0_mxn2v0x1_2_zn mux_0_mxn2v0x1_1_w_n4_32# 9.3fF
C120 totdiff3_1_diff2_0_an2v0x2_1_a totdiff3_1_diff2_0_in_b 2.0fF
C121 mux_0_gnd comp_0_an2v0x2_1_z 8.7fF
C122 totdiff3_1_mux_0_b0 totdiff3_1_mux_0_mxn2v0x1_0_zn 2.7fF
C123 totdiff3_1_diff2_2_an2v0x2_1_zn mux_0_vdd 8.8fF
C124 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_a0 4.8fF
C125 totdiff3_1_diff2_0_an2v0x2_2_zn mux_0_vdd 10.3fF
C126 mux_0_vdd totdiff3_1_mux_0_a1 38.7fF
C127 comp_0_an3v0x2_3_zn mux_0_gnd 8.8fF
C128 totdiff3_1_diff2_0_xnr2v8x05_0_zn mux_0_gnd 15.0fF
C129 totdiff3_1_diff2_2_xor3v1x2_0_cn mux_0_vdd 31.6fF
C130 totdiff3_0_mux_0_a2 mux_0_vdd 36.7fF
C131 totdiff3_0_diff2_0_xor3v1x2_0_cn mux_0_gnd 19.1fF
C132 totdiff3_0_diff2_2_xnr2v8x05_0_bn mux_0_gnd 6.7fF
C133 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# mux_0_b1 2.3fF
C134 totdiff3_0_diff2_0_an2v0x2_1_a totdiff3_0_diff2_0_in_b 2.0fF
C135 comp_0_nd3v0x2_0_a mux_0_vdd 9.6fF
C136 totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# 15.2fF
C137 mux_0_a0 mux_0_vdd 43.3fF
C138 mux_0_vdd totdiff3_1_diff2_0_xor3v1x2_0_cn 31.6fF
C139 totdiff3_1_diff2_2_in_a mux_0_gnd 27.8fF
C140 mux_0_a1 mux_0_mxn2v0x1_1_w_n4_32# 13.4fF
C141 comp_0_an3v0x2_0_zn mux_0_gnd 8.8fF
C142 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_0_mux_0_a0 4.8fF
C143 totdiff3_0_diff2_1_an2v0x2_1_zn mux_0_vdd 8.8fF
C144 totdiff3_0_diff2_2_in_b mux_0_gnd 60.5fF
C145 comp_0_an3v0x2_2_w_n4_32# comp_0_nd3v0x2_0_a 6.2fF
C146 totdiff3_0_diff2_0_xor3v1x2_0_cn totdiff3_0_diff2_0_xor3v1x2_0_zn 4.5fF
C147 mux_0_gnd totdiff3_1_diff2_1_an2v0x2_1_z 10.2fF
C148 mux_0_gnd mux_0_b0 9.4fF
C149 mux_0_gnd totdiff3_1_diff2_0_xor2v2x2_0_bn 11.2fF
C150 totdiff3_1_diff2_2_xor2v2x2_0_an mux_0_gnd 21.6fF
C151 comp_0_an3v0x2_2_w_n4_32# mux_0_a0 8.7fF
C152 totdiff3_0_diff2_0_an2v0x2_2_a mux_0_gnd 25.9fF
C153 totdiff3_1_diff2_0_or2v0x3_0_zn mux_0_gnd 9.0fF
C154 totdiff3_0_diff2_1_an2v0x2_2_zn mux_0_gnd 8.9fF
C155 mux_0_vdd totdiff3_1_diff2_0_an2v0x2_0_b 20.5fF
C156 totdiff3_0_diff2_0_xor3v1x2_0_iz mux_0_vdd 15.8fF
C157 totdiff3_0_diff2_2_xor2v2x2_0_an mux_0_vdd 25.5fF
C158 mux_0_vdd totdiff3_1_diff2_0_xor3v1x2_0_bn 15.4fF
C159 mux_0_b0 totdiff3_1_mux_0_a0 2.3fF
C160 totdiff3_0_diff2_2_in_a totdiff3_0_diff2_2_an2v0x2_0_zn 2.2fF
C161 mux_0_gnd totdiff3_1_mux_0_b0 10.9fF
C162 totdiff3_0_diff2_2_or2v0x3_0_zn mux_0_vdd 12.7fF
C163 totdiff3_1_mux_0_b1 mux_0_vdd 13.1fF
C164 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# mux_0_vdd 59.4fF
C165 mux_0_mxn2v0x1_0_w_n4_32# mux_0_a0 11.6fF
C166 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_b1 6.6fF
C167 totdiff3_0_mux_0_mxn2v0x1_2_zn totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# 8.9fF
C168 mux_0_mxn2v0x1_2_w_n4_n4# mux_0_o2 2.3fF
C169 totdiff3_0_diff2_1_in_c mux_0_gnd 34.1fF
C170 mux_0_mxn2v0x1_1_w_n4_32# mux_0_o2 6.3fF
C171 totdiff3_0_diff2_0_an2v0x2_1_z mux_0_vdd 17.9fF
C172 totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_xor3v1x2_0_cn 4.1fF
C173 totdiff3_1_diff2_2_xor3v1x2_0_bn mux_0_vdd 15.4fF
C174 mux_0_mxn2v0x1_1_w_n4_32# mux_0_b1 6.6fF
C175 comp_0_an3v0x2_0_z mux_0_vdd 2.3fF
C176 mux_0_vdd totdiff3_1_diff2_1_xor3v1x2_0_bn 15.4fF
C177 totdiff3_1_diff2_0_xor3v1x2_0_zn totdiff3_1_diff2_0_in_b 4.3fF
C178 totdiff3_0_diff2_2_an2v0x2_1_a mux_0_vdd 12.4fF
C179 totdiff3_1_diff2_2_in_c mux_0_vdd 40.7fF
C180 totdiff3_0_diff2_0_xor3v1x2_0_bn mux_0_gnd 9.1fF
C181 totdiff3_0_diff2_2_xnr2v8x05_0_an mux_0_gnd 5.5fF
C182 mux_0_a1 mux_0_gnd 33.3fF
C183 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_1_mux_0_mxn2v0x1_2_sn 9.2fF
C184 totdiff3_1_diff2_0_an2v0x2_1_a mux_0_gnd 20.0fF
C185 comp_0_an2v0x2_0_zn mux_0_gnd 8.9fF
C186 mux_0_vdd totdiff3_1_diff2_1_an2v0x2_2_a 59.6fF
C187 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_1_mux_0_a1 13.4fF
C188 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_xor3v1x2_0_cn 4.5fF
C189 comp_0_an2v0x2_3_b mux_0_gnd 15.0fF
C190 totdiff3_0_mux_0_b1 mux_0_vdd 13.1fF
C191 comp_0_an3v0x2_2_w_n4_32# comp_0_an3v0x2_0_z 9.5fF
C192 totdiff3_1_diff2_2_xor2v2x2_0_bn mux_0_gnd 11.2fF
C193 mux_0_mxn2v0x1_2_w_n4_n4# mux_0_mxn2v0x1_2_sn 9.2fF
C194 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_1_mux_0_mxn2v0x1_2_sn 9.3fF
C195 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_mxn2v0x1_1_zn 8.9fF
C196 mux_0_mxn2v0x1_2_sn mux_0_mxn2v0x1_1_w_n4_32# 9.3fF
C197 comp_0_nd3v0x2_0_c mux_0_gnd 18.9fF
C198 totdiff3_0_diff2_1_an2v0x2_2_a mux_0_vdd 59.6fF
C199 comp_0_an2v0x2_4_z mux_0_vdd 10.7fF
C200 totdiff3_0_diff2_2_xor3v1x2_0_iz mux_0_gnd 24.9fF
C201 totdiff3_0_diff2_1_an2v0x2_0_zn totdiff3_0_diff2_1_in_a 2.2fF
C202 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_mux_0_a2 4.1fF
C203 comp_0_an3v0x2_3_z mux_0_gnd 10.6fF
C204 comp_0_an3v0x2_2_z mux_0_gnd 10.7fF
C205 comp_0_an3v0x2_2_w_n4_32# mux_0_vdd 88.5fF
C206 totdiff3_0_mux_0_s totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 30.3fF
C207 mux_0_gnd totdiff3_1_diff2_0_xnr2v8x05_0_bn 7.5fF
C208 mux_0_mxn2v0x1_2_w_n4_n4# mux_0_s 15.2fF
C209 totdiff3_1_diff2_1_xnr2v8x05_0_an mux_0_gnd 5.5fF
C210 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_mux_0_a1 4.6fF
C211 mux_0_s mux_0_mxn2v0x1_1_w_n4_32# 36.4fF
C212 totdiff3_1_diff2_1_an2v0x2_1_a totdiff3_1_diff2_1_in_b 2.0fF
C213 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_1_mux_0_a1 4.8fF
C214 comp_0_an2v0x2_1_zn mux_0_gnd 8.9fF
C215 totdiff3_0_diff2_0_an2v0x2_2_zn mux_0_gnd 8.9fF
C216 totdiff3_0_diff2_1_xor3v1x2_0_iz mux_0_vdd 15.8fF
C217 mux_0_gnd totdiff3_1_mux_0_b2 11.9fF
C218 totdiff3_0_diff2_2_in_a mux_0_gnd 27.8fF
C219 totdiff3_1_diff2_2_xnr2v8x05_0_bn mux_0_vdd 14.4fF
C220 mux_0_mxn2v0x1_0_w_n4_32# mux_0_vdd 22.4fF
C221 totdiff3_0_diff2_2_an2v0x2_1_z mux_0_vdd 17.9fF
C222 mux_0_gnd mux_0_b1 12.7fF
C223 mux_0_gnd totdiff3_1_diff2_1_xor3v1x2_0_iz 24.9fF
C224 totdiff3_0_diff2_1_xor2v2x2_0_bn mux_0_vdd 17.7fF
C225 totdiff3_0_diff2_1_in_2c mux_0_vdd 34.0fF
C226 comp_0_nr3v0x2_0_z mux_0_vdd 8.7fF
C227 mux_0_vdd totdiff3_1_diff2_0_in_a 24.6fF
C228 totdiff3_0_mux_0_b1 totdiff3_0_diff2_1_xor2v2x2_0_bn 2.7fF
C229 mux_0_gnd totdiff3_1_diff2_0_an2v0x2_1_z 10.2fF
C230 totdiff3_1_diff2_2_an2v0x2_0_zn mux_0_gnd 8.9fF
C231 totdiff3_1_mux_0_b1 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 6.6fF
C232 mux_0_gnd totdiff3_1_diff2_0_an2v0x2_0_z 12.8fF
C233 totdiff3_0_mux_0_a0 totdiff3_0_diff2_0_xor3v1x2_0_cn 4.1fF
C234 totdiff3_1_mux_0_a2 mux_0_vdd 36.7fF
C235 totdiff3_0_diff2_1_an2v0x2_1_a mux_0_vdd 12.4fF
C236 comp_0_an3v0x2_2_w_n4_32# comp_0_nr3v0x2_0_z 21.8fF
C237 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# mux_0_a2 6.3fF
C238 totdiff3_1_diff2_2_an2v0x2_0_b mux_0_vdd 20.5fF
C239 mux_0_vdd totdiff3_1_diff2_1_in_c 39.6fF
C240 totdiff3_1_mux_0_mxn2v0x1_2_zn totdiff3_1_mux_0_b2 2.7fF
C241 mux_0_vdd totdiff3_1_diff2_1_in_a 24.6fF
C242 totdiff3_1_diff2_2_xnr2v8x05_0_an mux_0_gnd 5.5fF
C243 totdiff3_1_diff2_1_an2v0x2_0_b mux_0_vdd 20.5fF
C244 mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_zn 13.9fF
C245 comp_0_nd3v0x2_0_z mux_0_vdd 6.1fF
C246 totdiff3_1_diff2_2_in_2c mux_0_gnd 17.8fF
C247 totdiff3_1_mux_0_b1 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# 10.2fF
C248 totdiff3_0_diff2_2_an2v0x2_0_b mux_0_vdd 20.5fF
C249 mux_0_s mux_0_gnd 4.9fF
C250 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# mux_0_vdd 59.4fF
C251 mux_0_gnd totdiff3_1_diff2_0_xnr2v8x05_0_an 6.8fF
C252 totdiff3_0_diff2_2_xor3v1x2_0_zn totdiff3_0_mux_0_a2 4.6fF
C253 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_0_mux_0_mxn2v0x1_0_zn 8.9fF
C254 mux_0_a2 mux_0_vdd 27.5fF
C255 totdiff3_1_diff2_1_an2v0x2_1_a mux_0_gnd 20.0fF
C256 totdiff3_0_diff2_2_xor3v1x2_0_cn mux_0_vdd 31.6fF
C257 totdiff3_1_diff2_2_an2v0x2_2_zn mux_0_vdd 8.8fF
C258 totdiff3_0_diff2_0_xnr2v8x05_0_zn mux_0_vdd 4.4fF
C259 totdiff3_0_diff2_1_or2v0x3_0_zn mux_0_vdd 12.7fF
C260 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# mux_0_a0 5.1fF
C261 comp_0_an3v0x2_2_w_n4_32# comp_0_nd3v0x2_0_z 5.2fF
C262 totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_xor3v1x2_0_zn 4.6fF
C263 totdiff3_1_diff2_0_xor3v1x2_0_bn totdiff3_1_diff2_0_in_b 2.6fF
C264 totdiff3_0_mux_0_mxn2v0x1_0_sn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# 9.3fF
C265 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_0_mux_0_a1 4.8fF
C266 mux_0_o0 mux_0_a0 2.3fF
C267 comp_0_an3v0x2_2_w_n4_32# mux_0_a2 12.2fF
C268 comp_0_an3v0x2_1_a comp_0_or3v0x2_0_zn 4.1fF
C269 mux_0_a0 comp_0_an2v0x2_0_b 4.9fF
C270 totdiff3_0_diff2_2_xor3v1x2_0_bn totdiff3_0_diff2_2_in_b 2.6fF
C271 mux_0_gnd totdiff3_1_diff2_0_xor2v2x2_0_an 21.6fF
C272 comp_0_an2v0x2_3_z mux_0_gnd 20.8fF
C273 totdiff3_0_diff2_1_xnr2v8x05_0_zn totdiff3_0_diff2_1_in_c 3.1fF
C274 totdiff3_1_diff2_2_an2v0x2_1_a mux_0_gnd 20.0fF
C275 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_1_mux_0_mxn2v0x1_0_sn 9.2fF
C276 comp_0_nr2v0x2_1_a comp_0_nd3v0x2_0_c 3.8fF
C277 totdiff3_0_diff2_1_xnr2v8x05_0_bn mux_0_vdd 14.4fF
C278 totdiff3_0_diff2_1_an2v0x2_0_b mux_0_vdd 20.5fF
C279 totdiff3_1_diff2_2_in_b mux_0_gnd 60.5fF
C280 totdiff3_1_mux_0_a2 totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# 4.8fF
C281 mux_0_vdd totdiff3_1_diff2_0_in_b 50.3fF
C282 totdiff3_1_diff2_2_an2v0x2_1_zn mux_0_gnd 8.9fF
C283 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_1_mux_0_s 18.7fF
C284 mux_0_gnd totdiff3_1_diff2_0_an2v0x2_2_zn 8.9fF
C285 mux_0_gnd totdiff3_1_mux_0_a1 15.3fF
C286 totdiff3_1_diff2_1_xor3v1x2_0_bn totdiff3_1_diff2_1_in_b 2.6fF
C287 totdiff3_1_diff2_2_xor3v1x2_0_cn mux_0_gnd 18.8fF
C288 totdiff3_1_mux_0_a2 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 11.6fF
C289 totdiff3_0_mux_0_a2 mux_0_gnd 14.9fF
C290 totdiff3_1_diff2_2_in_c totdiff3_1_diff2_2_xnr2v8x05_0_zn 3.1fF
C291 mux_0_o0 mux_0_mxn2v0x1_0_w_n4_n4# 2.3fF
C292 totdiff3_1_diff2_2_xnr2v8x05_0_zn mux_0_vdd 4.4fF
C293 comp_0_nd3v0x2_0_a mux_0_gnd 21.1fF
C294 totdiff3_0_diff2_0_xnr2v8x05_0_bn mux_0_vdd 14.4fF
C295 mux_0_vdd totdiff3_1_diff2_1_in_b 50.3fF
C296 totdiff3_1_diff2_2_xor3v1x2_0_iz totdiff3_1_diff2_2_xor3v1x2_0_bn 2.4fF
C297 totdiff3_0_diff2_2_an2v0x2_1_zn mux_0_vdd 8.8fF
C298 totdiff3_0_diff2_2_an2v0x2_0_zn mux_0_vdd 8.8fF
C299 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# mux_0_vdd 20.7fF
C300 mux_0_gnd mux_0_a0 62.5fF
C301 mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_cn 19.1fF
C302 comp_0_an3v0x2_1_a comp_0_an3v0x2_0_zn 2.5fF
C303 totdiff3_0_diff2_1_an2v0x2_1_zn mux_0_gnd 8.9fF
C304 mux_0_mxn2v0x1_1_w_n4_32# mux_0_vdd 59.4fF
C305 totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_xor3v1x2_0_zn 4.6fF
C306 totdiff3_0_diff2_2_xor3v1x2_0_zn mux_0_vdd 18.9fF
C307 totdiff3_1_diff2_2_xor3v1x2_0_iz mux_0_vdd 15.8fF
C308 totdiff3_0_diff2_1_an2v0x2_0_z mux_0_vdd 24.6fF
C309 totdiff3_0_mux_0_b0 mux_0_vdd 28.1fF
C310 totdiff3_0_mux_0_b1 totdiff3_0_mux_0_b0 18.4fF
C311 totdiff3_0_mux_0_mxn2v0x1_2_sn totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# 9.2fF
C312 comp_0_an2v0x2_0_b mux_0_vdd 49.9fF
C313 totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_mux_0_a1 4.1fF
C314 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_o1 2.3fF
C315 totdiff3_1_mux_0_a0 totdiff3_1_diff2_0_xor3v1x2_0_cn 4.1fF
C316 mux_0_a0 comp_0_an2v0x2_1_b 2.2fF
C317 mux_0_gnd totdiff3_1_diff2_0_an2v0x2_0_b 7.3fF
C318 totdiff3_0_diff2_2_xor3v1x2_0_bn totdiff3_0_diff2_2_xor3v1x2_0_iz 2.4fF
C319 totdiff3_0_diff2_0_xor3v1x2_0_iz mux_0_gnd 25.5fF
C320 totdiff3_0_diff2_2_an2v0x2_2_z mux_0_vdd 2.4fF
C321 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_0_mux_0_mxn2v0x1_1_sn 9.2fF
C322 totdiff3_0_diff2_2_xor2v2x2_0_an mux_0_gnd 21.6fF
C323 mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_bn 9.1fF
C324 mux_0_mxn2v0x1_1_sn mux_0_mxn2v0x1_0_w_n4_n4# 9.2fF
C325 totdiff3_0_diff2_2_or2v0x3_0_zn mux_0_gnd 9.0fF
C326 totdiff3_1_mux_0_b1 mux_0_gnd 17.2fF
C327 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# mux_0_b0 5.2fF
C328 mux_0_mxn2v0x1_1_w_n4_32# mux_0_mxn2v0x1_1_zn 9.3fF
C329 totdiff3_0_diff2_0_xor3v1x2_0_bn totdiff3_0_diff2_0_in_b 2.6fF
C330 mux_0_a1 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 2.3fF
C331 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_gnd 80.2fF
C332 totdiff3_0_diff2_0_an2v0x2_1_z mux_0_gnd 10.2fF
C333 mux_0_o0 mux_0_mxn2v0x1_0_w_n4_32# 5.0fF
C334 totdiff3_1_mux_0_b1 totdiff3_1_diff2_1_xor2v2x2_0_bn 2.7fF
C335 mux_0_gnd totdiff3_1_diff2_2_xor3v1x2_0_bn 9.1fF
C336 totdiff3_0_diff2_0_xor2v2x2_0_bn mux_0_vdd 18.7fF
C337 comp_0_an3v0x2_0_z mux_0_gnd 36.9fF
C338 mux_0_gnd totdiff3_1_diff2_1_xor3v1x2_0_bn 9.1fF
C339 totdiff3_0_diff2_2_an2v0x2_1_a mux_0_gnd 20.0fF
C340 totdiff3_0_diff2_1_in_b mux_0_vdd 50.3fF
C341 totdiff3_1_diff2_2_in_c mux_0_gnd 35.0fF
C342 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_1_mux_0_b0 6.6fF
C343 totdiff3_1_diff2_0_an2v0x2_1_zn mux_0_vdd 8.8fF
C344 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_mux_0_b2 3.9fF
C345 totdiff3_0_diff2_1_xnr2v8x05_0_an mux_0_vdd 9.9fF
C346 mux_0_gnd mux_0_vdd 92.6fF
C347 mux_0_gnd totdiff3_1_diff2_1_an2v0x2_2_a 25.9fF
C348 totdiff3_0_mux_0_b1 mux_0_gnd 17.2fF
C349 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_b2 6.6fF
C350 totdiff3_0_diff2_0_an2v0x2_1_zn mux_0_vdd 8.8fF
C351 totdiff3_1_diff2_1_xor2v2x2_0_bn mux_0_vdd 17.7fF
C352 comp_0_an2v0x2_4_z mux_0_gnd 9.8fF
C353 comp_0_or3v0x2_1_zn mux_0_vdd 9.0fF
C354 totdiff3_0_diff2_1_an2v0x2_2_a mux_0_gnd 25.9fF
C355 comp_0_an2v0x2_2_z mux_0_vdd 9.4fF
C356 comp_0_an2v0x2_3_zn mux_0_vdd 8.8fF
C357 totdiff3_1_diff2_0_xor3v1x2_0_iz totdiff3_1_diff2_0_xor3v1x2_0_bn 2.4fF
C358 totdiff3_0_diff2_1_xor3v1x2_0_bn mux_0_vdd 15.4fF
C359 totdiff3_1_diff2_2_xor3v1x2_0_cn totdiff3_1_diff2_2_an2v0x2_2_a 2.3fF
C360 totdiff3_0_diff2_0_xor3v1x2_0_zn mux_0_vdd 18.9fF
C361 mux_0_vdd totdiff3_1_mux_0_a0 35.4fF
C362 comp_0_an2v0x2_2_zn mux_0_vdd 8.8fF
C363 mux_0_vdd comp_0_an2v0x2_1_b 14.2fF
C364 mux_0_vdd totdiff3_1_diff2_1_xor3v1x2_0_zn 18.9fF
C365 totdiff3_1_mux_0_a1 totdiff3_1_diff2_1_xor3v1x2_0_cn 4.1fF
C366 totdiff3_0_diff2_2_xnr2v8x05_0_zn mux_0_vdd 4.4fF
C367 totdiff3_0_mux_0_b2 mux_0_vdd 3.1fF
C368 totdiff3_0_diff2_0_or2v0x3_0_zn mux_0_vdd 12.7fF
C369 totdiff3_0_diff2_1_xor3v1x2_0_iz mux_0_gnd 24.9fF
C370 mux_0_mxn2v0x1_2_w_n4_n4# mux_0_a2 4.8fF
C371 mux_0_mxn2v0x1_1_w_n4_32# mux_0_a2 11.6fF
C372 mux_0_mxn2v0x1_0_w_n4_32# mux_0_gnd 2.6fF
C373 totdiff3_1_diff2_2_xnr2v8x05_0_bn mux_0_gnd 6.7fF
C374 totdiff3_1_diff2_0_an2v0x2_0_zn mux_0_vdd 8.8fF
C375 totdiff3_0_diff2_0_in_a mux_0_vdd 24.6fF
C376 mux_0_vdd totdiff3_1_diff2_1_xnr2v8x05_0_zn 4.4fF
C377 totdiff3_0_diff2_2_xor3v1x2_0_cn totdiff3_0_diff2_2_xor3v1x2_0_zn 4.5fF
C378 totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# totdiff3_0_mux_0_a2 4.8fF
C379 totdiff3_0_diff2_2_an2v0x2_1_z mux_0_gnd 10.2fF
C380 mux_0_mxn2v0x1_0_zn mux_0_b0 2.7fF
C381 totdiff3_0_diff2_2_xor2v2x2_0_an totdiff3_0_diff2_2_xor2v2x2_0_bn 3.3fF
C382 mux_0_mxn2v0x1_2_zn mux_0_b2 2.7fF
C383 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_1_mux_0_mxn2v0x1_0_zn 8.9fF
C384 mux_0_vdd totdiff3_1_diff2_0_xor3v1x2_0_iz 15.8fF
C385 totdiff3_0_diff2_1_xor3v1x2_0_iz totdiff3_0_diff2_1_xor3v1x2_0_bn 2.4fF
C386 totdiff3_0_diff2_1_in_2c mux_0_gnd 17.5fF
C387 totdiff3_0_diff2_1_xor2v2x2_0_bn mux_0_gnd 11.2fF
C388 comp_0_an3v0x2_2_b mux_0_vdd 39.7fF
C389 comp_0_nr3v0x2_0_z mux_0_gnd 21.2fF
C390 totdiff3_0_diff2_0_an2v0x2_0_z mux_0_vdd 24.6fF
C391 mux_0_gnd totdiff3_1_diff2_0_in_a 28.0fF
C392 comp_0_an2v0x2_4_zn mux_0_vdd 8.8fF
C393 totdiff3_0_diff2_1_in_b totdiff3_0_diff2_1_an2v0x2_1_a 2.0fF
C394 comp_0_an3v0x2_1_zn mux_0_vdd 4.9fF
C395 totdiff3_0_diff2_0_an2v0x2_2_a totdiff3_0_diff2_0_xor3v1x2_0_cn 2.3fF
C396 totdiff3_1_diff2_2_or2v0x3_0_zn mux_0_vdd 12.7fF
C397 totdiff3_1_mux_0_a2 mux_0_gnd 14.9fF
C398 totdiff3_0_diff2_1_an2v0x2_1_a mux_0_gnd 20.0fF
C399 totdiff3_0_diff2_2_in_c mux_0_vdd 40.7fF
C400 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_0_mux_0_mxn2v0x1_1_zn 8.9fF
C401 comp_0_an3v0x2_2_w_n4_32# comp_0_an3v0x2_2_b 21.4fF
C402 mux_0_gnd totdiff3_1_diff2_2_an2v0x2_0_b 5.9fF
C403 totdiff3_0_diff2_0_xor2v2x2_0_an mux_0_vdd 27.4fF
C404 mux_0_gnd totdiff3_1_diff2_1_in_c 34.1fF
C405 mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# 26.1fF
C406 totdiff3_0_mux_0_a0 mux_0_a0 2.3fF
C407 mux_0_gnd totdiff3_1_diff2_1_in_a 27.8fF
C408 comp_0_an3v0x2_1_zn comp_0_an3v0x2_2_w_n4_32# 5.8fF
C409 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_in_b 4.3fF
C410 totdiff3_1_diff2_1_an2v0x2_0_b mux_0_gnd 5.9fF
C411 totdiff3_0_diff2_2_xor2v2x2_0_bn mux_0_vdd 17.7fF
C412 totdiff3_1_mux_0_b1 totdiff3_1_diff2_1_xor2v2x2_0_an 3.9fF
C413 comp_0_nd3v0x2_0_z mux_0_gnd 5.3fF
C414 totdiff3_1_diff2_1_in_2c mux_0_vdd 34.0fF
C415 totdiff3_0_diff2_2_an2v0x2_0_b mux_0_gnd 5.9fF
C416 totdiff3_1_diff2_0_an2v0x2_0_zn totdiff3_1_diff2_0_in_a 2.2fF
C417 totdiff3_0_diff2_2_an2v0x2_2_a mux_0_vdd 59.6fF
C418 mux_0_a1 comp_0_an3v0x2_3_zn 3.6fF
C419 mux_0_a2 mux_0_gnd 35.4fF
C420 totdiff3_0_diff2_0_an2v0x2_0_b mux_0_vdd 20.5fF
C421 totdiff3_0_diff2_2_xor3v1x2_0_cn mux_0_gnd 18.8fF
C422 mux_0_gnd totdiff3_1_diff2_2_an2v0x2_2_zn 8.9fF
C423 totdiff3_1_diff2_2_an2v0x2_2_z mux_0_vdd 2.4fF
C424 totdiff3_0_diff2_0_xnr2v8x05_0_zn mux_0_gnd 15.0fF
C425 totdiff3_0_diff2_1_or2v0x3_0_zn mux_0_gnd 9.0fF
C426 totdiff3_1_mux_0_b0 totdiff3_1_diff2_0_xor2v2x2_0_bn 2.7fF
C427 mux_0_vdd totdiff3_1_diff2_2_an2v0x2_2_a 59.6fF
C428 totdiff3_1_diff2_2_xor3v1x2_0_zn totdiff3_1_diff2_2_xor3v1x2_0_cn 4.5fF
C429 totdiff3_1_diff2_1_an2v0x2_0_z mux_0_vdd 24.6fF
C430 mux_0_vdd totdiff3_1_diff2_1_xor2v2x2_0_an 25.5fF
C431 totdiff3_0_mux_0_b0 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# 6.6fF
C432 mux_0_gnd totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# 76.2fF
C433 comp_0_nr2v0x2_1_a mux_0_vdd 7.1fF
C434 totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_1_mux_0_mxn2v0x1_1_sn 9.3fF
C435 totdiff3_1_mux_0_mxn2v0x1_2_zn totdiff3_1_mux_0_mxn2v0x1_2_w_n4_n4# 8.9fF
C436 totdiff3_1_diff2_1_an2v0x2_2_zn mux_0_vdd 8.8fF
C437 totdiff3_1_diff2_1_in_c totdiff3_1_diff2_1_xnr2v8x05_0_zn 3.1fF
C438 mux_0_vdd totdiff3_1_diff2_1_xor3v1x2_0_cn 31.6fF
C439 totdiff3_1_diff2_1_an2v0x2_2_a totdiff3_1_diff2_1_xor3v1x2_0_cn 2.3fF
C440 totdiff3_1_diff2_1_an2v0x2_1_zn mux_0_vdd 8.8fF
C441 totdiff3_0_diff2_1_xor3v1x2_0_zn mux_0_vdd 18.9fF
C442 totdiff3_0_diff2_1_xnr2v8x05_0_bn mux_0_gnd 6.7fF
C443 totdiff3_0_diff2_1_an2v0x2_0_b mux_0_gnd 5.9fF
C444 totdiff3_1_mux_0_mxn2v0x1_2_zn totdiff3_1_mux_0_mxn2v0x1_1_w_n4_32# 9.3fF
C445 totdiff3_0_diff2_0_an2v0x2_1_a mux_0_vdd 12.4fF
C446 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_mxn2v0x1_0_sn 9.2fF
C447 comp_0_nr3v0x2_0_a mux_0_vdd 4.0fF
C448 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_1_mux_0_a0 4.8fF
C449 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_diff2_2_xor2v2x2_0_bn 3.3fF
C450 totdiff3_0_diff2_1_in_a mux_0_vdd 24.6fF
C451 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_n4# totdiff3_1_mux_0_mxn2v0x1_1_sn 9.2fF
C452 totdiff3_0_mux_0_s totdiff3_0_mux_0_a2 4.5fF
C453 totdiff3_0_mux_0_a0 mux_0_vdd 35.4fF
C454 mux_0_gnd totdiff3_1_diff2_0_in_b 60.8fF
C455 totdiff3_0_diff2_1_xnr2v8x05_0_zn mux_0_vdd 4.4fF
C456 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# mux_0_a0 2.3fF
C457 totdiff3_0_diff2_1_an2v0x2_1_z mux_0_vdd 17.9fF
C458 comp_0_an3v0x2_2_w_n4_32# comp_0_nr3v0x2_0_a 15.0fF
C459 mux_0_mxn2v0x1_1_w_n4_32# mux_0_o1 5.0fF
C460 totdiff3_0_diff2_1_xor2v2x2_0_an mux_0_vdd 25.5fF
C461 totdiff3_1_diff2_1_or2v0x3_0_zn mux_0_vdd 12.7fF
C462 totdiff3_0_mux_0_b1 totdiff3_0_diff2_1_xor2v2x2_0_an 3.9fF
C463 totdiff3_0_mux_0_mxn2v0x1_0_sn totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 9.2fF
C464 mux_0_gnd totdiff3_1_diff2_2_xnr2v8x05_0_zn 11.9fF
C465 totdiff3_0_diff2_0_xnr2v8x05_0_bn mux_0_gnd 7.5fF
C466 mux_0_gnd totdiff3_1_diff2_1_in_b 60.5fF
C467 mux_0_mxn2v0x1_1_sn mux_0_mxn2v0x1_1_w_n4_32# 9.3fF
C468 totdiff3_0_mux_0_b0 totdiff3_0_diff2_0_xor2v2x2_0_bn 2.7fF
C469 totdiff3_0_diff2_2_an2v0x2_1_zn mux_0_gnd 8.9fF
C470 totdiff3_1_diff2_2_xor2v2x2_0_an totdiff3_1_mux_0_b2 3.9fF
C471 totdiff3_0_diff2_2_an2v0x2_0_zn mux_0_gnd 8.9fF
C472 comp_0_an3v0x2_1_a mux_0_a0 6.8fF
C473 mux_0_mxn2v0x1_2_w_n4_n4# mux_0_gnd 25.5fF
C474 totdiff3_0_diff2_0_xnr2v8x05_0_an mux_0_vdd 9.9fF
C475 totdiff3_1_diff2_0_an2v0x2_2_a totdiff3_1_diff2_0_xor3v1x2_0_cn 2.3fF
C476 comp_0_an3v0x2_2_zn mux_0_vdd 4.9fF
C477 totdiff3_0_diff2_2_xor3v1x2_0_zn mux_0_gnd 11.9fF
C478 totdiff3_1_diff2_2_in_a totdiff3_1_diff2_2_an2v0x2_0_zn 2.2fF
C479 totdiff3_1_diff2_2_xor3v1x2_0_iz mux_0_gnd 24.9fF
C480 totdiff3_0_mux_0_b0 mux_0_gnd 10.9fF
C481 totdiff3_0_diff2_1_an2v0x2_0_z mux_0_gnd 12.8fF
C482 totdiff3_0_diff2_2_xor3v1x2_0_bn mux_0_vdd 15.4fF
C483 totdiff3_0_diff2_2_an2v0x2_2_zn mux_0_vdd 8.8fF
C484 totdiff3_1_diff2_2_xor3v1x2_0_zn mux_0_vdd 18.9fF
C485 mux_0_gnd comp_0_an2v0x2_0_b 32.8fF
C486 totdiff3_1_diff2_1_xor3v1x2_0_zn totdiff3_1_diff2_1_in_b 4.3fF
C487 comp_0_an3v0x2_2_zn comp_0_an3v0x2_2_w_n4_32# 5.8fF
C488 totdiff3_0_diff2_2_an2v0x2_2_a totdiff3_0_diff2_2_xor3v1x2_0_cn 2.3fF
C489 mux_0_mxn2v0x1_0_sn mux_0_mxn2v0x1_0_w_n4_32# 9.3fF
C490 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_s 36.4fF
C491 mux_0_vdd totdiff3_1_diff2_1_xnr2v8x05_0_bn 14.4fF
C492 totdiff3_0_diff2_2_an2v0x2_2_z mux_0_gnd 2.5fF
C493 totdiff3_0_diff2_1_xor2v2x2_0_bn totdiff3_0_diff2_1_xor2v2x2_0_an 3.3fF
C494 totdiff3_0_diff2_2_an2v0x2_0_z mux_0_vdd 24.6fF
C495 totdiff3_0_diff2_0_in_b mux_0_vdd 50.3fF
C496 totdiff3_0_mux_0_b1 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_n4# 10.2fF
C497 totdiff3_0_diff2_0_xor2v2x2_0_bn mux_0_gnd 11.2fF
C498 totdiff3_0_mux_0_s mux_0_vdd 7.9fF
C499 totdiff3_1_diff2_2_xor2v2x2_0_bn totdiff3_1_mux_0_b2 2.7fF
C500 totdiff3_0_diff2_1_in_b mux_0_gnd 60.5fF
C501 totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# mux_0_a2 2.3fF
C502 totdiff3_1_diff2_0_an2v0x2_1_zn mux_0_gnd 8.9fF
C503 comp_0_nr3v0x2_0_a mux_0_a2 2.5fF
C504 totdiff3_0_diff2_1_xnr2v8x05_0_an mux_0_gnd 5.5fF
C505 comp_0_an3v0x2_1_a mux_0_vdd 72.4fF
C506 mux_0_a0 comp_0_or3v0x2_0_zn 3.3fF
C507 mux_0_vdd totdiff3_1_diff2_0_an2v0x2_2_a 61.1fF
C508 totdiff3_0_diff2_0_an2v0x2_1_zn mux_0_gnd 8.9fF
C509 comp_0_an3v0x2_2_b comp_0_an2v0x2_0_b 2.5fF
C510 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_mxn2v0x1_2_zn 9.3fF
C511 totdiff3_1_diff2_1_an2v0x2_0_zn mux_0_vdd 8.8fF
C512 totdiff3_0_diff2_1_xor3v1x2_0_bn totdiff3_0_diff2_1_in_b 2.6fF
C513 mux_0_gnd totdiff3_1_diff2_1_xor2v2x2_0_bn 11.2fF
C514 comp_0_an2v0x2_2_z mux_0_gnd 11.1fF
C515 comp_0_or3v0x2_1_zn mux_0_gnd 10.9fF
C516 mux_0_gnd comp_0_an2v0x2_3_zn 8.9fF
C517 totdiff3_1_diff2_0_xor2v2x2_0_bn totdiff3_1_diff2_0_xor2v2x2_0_an 3.3fF
C518 totdiff3_1_mux_0_a2 totdiff3_1_diff2_2_xor3v1x2_0_zn 4.6fF
C519 totdiff3_0_mux_0_b0 totdiff3_0_diff2_0_xor2v2x2_0_an 3.9fF
C520 totdiff3_0_diff2_1_xor3v1x2_0_bn mux_0_gnd 9.1fF
C521 comp_0_an3v0x2_2_w_n4_32# comp_0_an3v0x2_1_a 8.3fF
C522 totdiff3_0_diff2_0_xor3v1x2_0_zn mux_0_gnd 13.9fF
C523 mux_0_gnd totdiff3_1_mux_0_a0 14.9fF
C524 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# mux_0_vdd 21.4fF
C525 comp_0_an2v0x2_2_zn mux_0_gnd 8.9fF
C526 mux_0_gnd comp_0_an2v0x2_1_b 5.9fF
C527 mux_0_gnd totdiff3_1_diff2_1_xor3v1x2_0_zn 11.9fF
C528 totdiff3_0_diff2_2_xnr2v8x05_0_zn mux_0_gnd 11.9fF
C529 totdiff3_0_mux_0_b2 mux_0_gnd 11.9fF
C530 totdiff3_0_diff2_0_or2v0x3_0_zn mux_0_gnd 9.0fF
C531 totdiff3_0_diff2_0_an2v0x2_0_zn mux_0_vdd 8.8fF
C532 totdiff3_1_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_1_mux_0_mxn2v0x1_0_sn 9.3fF
C533 mux_0_gnd totdiff3_1_diff2_0_an2v0x2_0_zn 10.8fF
C534 totdiff3_0_diff2_0_in_a mux_0_gnd 28.0fF
C535 totdiff3_1_mux_0_b0 totdiff3_1_diff2_0_xor2v2x2_0_an 3.9fF
C536 mux_0_gnd totdiff3_1_diff2_1_xnr2v8x05_0_zn 11.9fF
C537 mux_0_vdd totdiff3_1_diff2_2_an2v0x2_0_z 24.6fF
C538 totdiff3_0_diff2_2_in_2c mux_0_vdd 33.2fF
C539 mux_0_gnd totdiff3_1_diff2_0_xor3v1x2_0_iz 25.5fF
C540 totdiff3_0_diff2_0_an2v0x2_0_z mux_0_gnd 12.8fF
C541 comp_0_an3v0x2_0_zn mux_0_a0 4.6fF
C542 mux_0_gnd comp_0_an3v0x2_2_b 23.0fF
C543 totdiff3_0_mux_0_mxn2v0x1_1_w_n4_32# totdiff3_0_mux_0_a1 13.4fF
C544 totdiff3_1_diff2_2_an2v0x2_1_z mux_0_vdd 17.9fF
C545 comp_0_an2v0x2_4_zn mux_0_gnd 8.9fF
C546 totdiff3_0_diff2_0_xor2v2x2_0_bn totdiff3_0_diff2_0_xor2v2x2_0_an 3.3fF
C547 comp_0_an3v0x2_1_zn mux_0_gnd 8.8fF
C548 totdiff3_0_diff2_1_xor3v1x2_0_cn mux_0_vdd 31.6fF
C549 totdiff3_0_diff2_1_an2v0x2_0_zn mux_0_vdd 8.8fF
C550 totdiff3_1_diff2_2_or2v0x3_0_zn mux_0_gnd 9.0fF
C551 totdiff3_0_diff2_2_in_c mux_0_gnd 35.0fF
C552 totdiff3_1_mux_0_s mux_0_vdd 7.9fF
C553 comp_0_or3v0x2_0_zn mux_0_vdd 9.0fF
C554 totdiff3_0_diff2_1_xor3v1x2_0_cn totdiff3_0_diff2_1_an2v0x2_2_a 2.3fF
C555 totdiff3_0_diff2_0_xor2v2x2_0_an mux_0_gnd 21.6fF
C556 totdiff3_0_mux_0_mxn2v0x1_0_w_n4_32# totdiff3_0_mux_0_a0 11.6fF
C557 mux_0_mxn2v0x1_0_zn mux_0_mxn2v0x1_0_w_n4_n4# 8.9fF
C558 totdiff3_0_diff2_2_xor2v2x2_0_bn mux_0_gnd 11.2fF
C559 totdiff3_0_mux_0_a1 mux_0_vdd 38.7fF
C560 mux_0_b2 mux_0_vdd 11.8fF
C561 totdiff3_1_diff2_1_an2v0x2_0_zn totdiff3_1_diff2_1_in_a 2.2fF
C562 totdiff3_0_mux_0_b1 totdiff3_0_mux_0_a1 39.4fF
C563 totdiff3_1_diff2_1_in_2c mux_0_gnd 17.5fF
C564 comp_0_an2v0x2_1_z mux_0_vdd 22.0fF
C565 totdiff3_0_diff2_2_an2v0x2_2_a mux_0_gnd 25.9fF
C566 totdiff3_0_diff2_2_in_c totdiff3_0_diff2_2_xnr2v8x05_0_zn 3.1fF
C567 mux_0_o0 mux_0_mxn2v0x1_0_sn 4.3fF
C568 comp_0_an3v0x2_3_zn mux_0_vdd 10.7fF
C569 totdiff3_0_diff2_0_an2v0x2_0_b mux_0_gnd 7.3fF
C570 totdiff3_1_diff2_0_xnr2v8x05_0_zn mux_0_vdd 4.4fF
C571 mux_0_gnd totdiff3_1_diff2_2_an2v0x2_2_z 2.5fF
C572 mux_0_gnd totdiff3_1_diff2_2_an2v0x2_2_a 25.9fF
C573 totdiff3_1_diff2_1_an2v0x2_0_z mux_0_gnd 12.8fF
C574 totdiff3_0_diff2_0_xor3v1x2_0_cn mux_0_vdd 31.6fF
C575 totdiff3_0_diff2_2_xnr2v8x05_0_bn mux_0_vdd 14.4fF
C576 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_b0 8.7fF
C577 mux_0_gnd totdiff3_1_diff2_1_xor2v2x2_0_an 21.6fF
C578 totdiff3_0_mux_0_b2 totdiff3_0_diff2_2_xor2v2x2_0_bn 2.7fF
C579 totdiff3_0_diff2_2_an2v0x2_1_a totdiff3_0_diff2_2_in_b 2.0fF
C580 comp_0_nr2v0x2_1_a mux_0_gnd 22.9fF
C581 totdiff3_1_diff2_1_an2v0x2_2_zn mux_0_gnd 8.9fF
C582 mux_0_gnd totdiff3_1_diff2_1_xor3v1x2_0_cn 18.8fF
C583 totdiff3_0_diff2_1_xor3v1x2_0_zn totdiff3_0_diff2_1_in_b 4.3fF
C584 totdiff3_1_diff2_2_in_a mux_0_vdd 24.6fF
C585 comp_0_an3v0x2_0_zn mux_0_vdd 10.7fF
C586 totdiff3_0_diff2_2_in_b mux_0_vdd 50.3fF
C587 totdiff3_1_diff2_1_xor2v2x2_0_bn totdiff3_1_diff2_1_xor2v2x2_0_an 3.3fF
C588 totdiff3_1_mux_0_b1 totdiff3_1_mux_0_b0 18.4fF
C589 mux_0_gnd totdiff3_1_diff2_1_an2v0x2_1_zn 8.9fF
C590 totdiff3_0_diff2_1_xor3v1x2_0_zn mux_0_gnd 11.9fF
C591 totdiff3_0_mux_0_mxn2v0x1_2_w_n4_n4# mux_0_gnd 25.5fF
C592 totdiff3_0_diff2_0_an2v0x2_1_a mux_0_gnd 20.0fF
C593 totdiff3_1_diff2_1_an2v0x2_1_z mux_0_vdd 17.9fF
C594 mux_0_vdd mux_0_b0 13.2fF
C595 mux_0_vdd totdiff3_1_diff2_0_xor2v2x2_0_bn 18.7fF
C596 totdiff3_1_mux_0_a2 totdiff3_1_mux_0_s 4.5fF
C597 totdiff3_1_diff2_2_xor2v2x2_0_an mux_0_vdd 25.5fF
C598 comp_0_nr3v0x2_0_a mux_0_gnd 19.9fF
C599 totdiff3_0_diff2_0_an2v0x2_2_a mux_0_vdd 61.1fF
C600 totdiff3_1_diff2_0_in_a 0 4.4fF
C601 totdiff3_1_diff2_0_an2v0x2_0_b 0 2.9fF
C602 totdiff3_1_diff2_1_in_c 0 37.1fF
C603 totdiff3_1_diff2_0_an2v0x2_0_z 0 5.0fF
C604 totdiff3_1_diff2_1_in_a 0 4.4fF
C605 totdiff3_1_mux_0_a1 0 28.9fF
C606 totdiff3_1_diff2_1_an2v0x2_0_b 0 2.9fF
C607 totdiff3_1_diff2_2_in_c 0 36.8fF
C608 totdiff3_1_diff2_1_an2v0x2_0_z 0 5.0fF
C609 totdiff3_1_diff2_1_in_2c 0 29.6fF
C610 totdiff3_1_diff2_2_in_a 0 4.4fF
C611 totdiff3_1_mux_0_a2 0 38.7fF
C612 totdiff3_1_diff2_2_an2v0x2_0_b 0 2.9fF
C613 totdiff3_1_diff2_2_an2v0x2_0_z 0 5.0fF
C614 totdiff3_1_diff2_2_in_2c 0 34.8fF
C615 totdiff3_1_mux_0_b0 0 47.5fF
C616 totdiff3_1_mux_0_s 0 16.3fF
C617 totdiff3_1_mux_0_a0 0 99.1fF
C618 totdiff3_1_mux_0_b1 0 87.1fF
C619 totdiff3_1_mux_0_b2 0 24.6fF
C620 mux_0_b2 0 43.5fF
C621 mux_0_b0 0 53.7fF
C622 mux_0_a1 0 43.2fF
C623 mux_0_a2 0 71.0fF
C624 mux_0_vdd 0 680.3fF
C625 mux_0_b1 0 32.9fF
C626 mux_0_a0 0 75.4fF
C627 mux_0_gnd 0 903.1fF
C628 comp_0_nr3v0x2_0_a 0 8.6fF
C629 totdiff3_0_diff2_0_in_a 0 4.4fF
C630 totdiff3_0_diff2_0_an2v0x2_0_b 0 2.9fF
C631 totdiff3_0_diff2_1_in_c 0 37.1fF
C632 totdiff3_0_diff2_0_an2v0x2_0_z 0 5.0fF
C633 totdiff3_0_diff2_1_in_a 0 4.4fF
C634 totdiff3_0_mux_0_a1 0 28.9fF
C635 totdiff3_0_diff2_1_an2v0x2_0_b 0 2.9fF
C636 totdiff3_0_diff2_2_in_c 0 36.8fF
C637 totdiff3_0_diff2_1_an2v0x2_0_z 0 5.0fF
C638 totdiff3_0_diff2_1_in_2c 0 29.6fF
C639 totdiff3_0_diff2_2_in_a 0 4.4fF
C640 totdiff3_0_mux_0_a2 0 38.7fF
C641 totdiff3_0_diff2_2_an2v0x2_0_b 0 2.9fF
C642 totdiff3_0_diff2_2_an2v0x2_0_z 0 5.0fF
C643 totdiff3_0_diff2_2_in_2c 0 34.8fF
C644 totdiff3_0_mux_0_b0 0 47.5fF
C645 totdiff3_0_mux_0_s 0 16.3fF
C646 totdiff3_0_mux_0_a0 0 99.1fF
C647 totdiff3_0_mux_0_b1 0 87.1fF
C648 totdiff3_0_mux_0_b2 0 24.6fF
C649 mux_0_s 0 9.4fF
C650 mux_0_o1 0 2.4fF

v_dd mux_0_vdd 0 5
v_ss mux_0_gnd 0 0

v_a11 totdiff3_0_diff2_0_in_a 0 DC 1 PULSE(5 0 0 0.1n 0.1n 15n 30n)
v_a12 totdiff3_0_diff2_1_in_a 0 DC 1 PULSE(5 0 0 0.1n 0.1n 15n 30n)
v_a13 totdiff3_0_diff2_2_in_a 0 DC 1 PULSE(5 0 0 0.1n 0.1n 15n 30n)
v_a21 totdiff3_1_diff2_0_in_a 0 DC 1 PULSE(5 0 0 0.1n 0.1n 15n 30n)
v_a22 totdiff3_1_diff2_1_in_a 0 DC 1 PULSE(5 0 0 0.1n 0.1n 15n 30n)
v_a23 totdiff3_1_diff2_2_in_a 0 DC 1 PULSE(5 0 0 0.1n 0.1n 15n 30n)

v_b11 totdiff3_0_diff2_0_in_b 0 DC 1 PULSE(5 0 0 0.1n 0.1n 30n 60n)
v_b12 totdiff3_0_diff2_1_in_b 0 DC 1 PULSE(5 0 0 0.1n 0.1n 30n 60n)
v_b13 totdiff3_0_diff2_2_in_b 0 DC 1 PULSE(5 0 0 0.1n 0.1n 30n 60n)
v_b21 totdiff3_1_diff2_0_in_b 0 DC 1 PULSE(5 0 0 0.1n 0.1n 30n 60n)
v_b22 totdiff3_1_diff2_1_in_b 0 DC 1 PULSE(5 0 0 0.1n 0.1n 30n 60n)
v_b23 totdiff3_1_diff2_2_in_b 0 DC 1 PULSE(5 0 0 0.1n 0.1n 30n 60n)
 
v_c2 mux_0_s 0  DC 1 PULSE(5 0 0 0.1n 0.1n 30n 60n)
.tran 0.1ns 200ns 

.control
run 
setplot tran1
plot comp_0_nd3v0x2_0_z
.endc 
