* Mon Aug 16 14:10:56 CEST 2004
.subckt an2v4x2 a b vdd vss z 
*SPICE circuit <an2v4x2> from XCircuit v3.10

m1 z n2 vdd vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m2 z n2 vss vss n w=14u l=2.3636u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m3 n1 a vss vss n w=7u l=2.3636u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m4 n2 a vdd vdd p w=8u l=2.3636u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
m5 n2 b n1 vss n w=7u l=2.3636u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m6 n2 b vdd vdd p w=8u l=2.3636u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
.ends
