* Sat Aug 27 22:10:21 CEST 2005
.subckt iv1v5x4 a vdd vss z 
*SPICE circuit <iv1v5x4> from XCircuit v3.20

m1 z a vss vss n w=22u l=2.3636u ad='22u*5u+12p' as='22u*5u+12p' pd='22u*2+14u' ps='22u*2+14u'
m2 z a vdd vdd p w=56u l=2.3636u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
.ends
