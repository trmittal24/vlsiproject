* Mon Aug 16 14:11:00 CEST 2004
.subckt nr3v0x2 a b c vdd vss z 
*SPICE circuit <nr3v0x2> from XCircuit v3.10

m1 z a vss vss n w=15u l=2u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m2 z c vss vss n w=15u l=2u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m3 n1 a vdd vdd p w=81u l=2u ad='81u*5u+12p' as='81u*5u+12p' pd='81u*2+14u' ps='81u*2+14u'
m4 n2 b n1 vdd p w=81u l=2u ad='81u*5u+12p' as='81u*5u+12p' pd='81u*2+14u' ps='81u*2+14u'
m5 z b vss vss n w=15u l=2u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m6 z c n2 vdd p w=81u l=2u ad='81u*5u+12p' as='81u*5u+12p' pd='81u*2+14u' ps='81u*2+14u'
.ends
