* Spice description of vfeed6
* Spice driver version 134999461
* Date 22/07/2007 at 11:00:26
* vsxlib 0.13um values
.subckt vfeed6 vdd vss
.ends
