* Spice description of or2v0x1
* Spice driver version 134999461
* Date 17/05/2007 at  9:32:38
* wsclib 0.13um values
.subckt or2v0x1 a b vdd vss z
M01 03    a     vdd   vdd p  L=0.12U  W=1.155U AS=0.306075P AD=0.306075P PS=2.84U   PD=2.84U
M02 sig1  a     vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M03 sig1  b     03    vdd p  L=0.12U  W=1.155U AS=0.306075P AD=0.306075P PS=2.84U   PD=2.84U
M04 vss   b     sig1  vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M5  vdd   sig1  z     vdd p  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
M6  vss   sig1  z     vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
C4  a     vss   0.367f
C5  b     vss   0.404f
C1  sig1  vss   0.592f
C3  z     vss   0.657f
.ends
