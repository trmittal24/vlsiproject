* Tue Apr  4 18:55:29 CEST 2006
.subckt iv1v8x1 a vdd vss z 
*SPICE circuit <iv1v8x1> from XCircuit v3.20

m1 z a vss vss n w=7u l=2.3636u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m2 z a vdd vdd p w=15u l=2.3636u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
.ends
