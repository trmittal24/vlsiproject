* Tue Apr  4 18:58:28 CEST 2006
.subckt iv1v3x3 a vdd vss z 
*SPICE circuit <iv1v3x3> from XCircuit v3.20

m1 z a vss vss n w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m2 z a vdd vdd p w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
.ends
