* Spice description of nr2v0x1
* Spice driver version 134999461
* Date 17/05/2007 at  9:25:34
* wsclib 0.13um values
.subckt nr2v0x1 a b vdd vss z
M01 vdd   a     01    vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M02 vss   a     z     vss n  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M03 01    b     z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M04 z     b     vss   vss n  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
C4  a     vss   0.287f
C3  b     vss   0.327f
C2  z     vss   0.745f
.ends
