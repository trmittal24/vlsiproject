magic
tech scmos
timestamp 1523171363
<< polysilicon >>
rect 1939 313 1941 324
rect 1868 246 1901 248
rect 1860 166 1903 168
rect 1967 85 1969 89
rect 1897 83 1969 85
rect 1897 64 1899 83
rect 1868 62 1899 64
rect 1903 -8 1905 9
rect 1925 -1 1927 8
rect 1925 -6 1927 -5
<< metal1 >>
rect 1930 328 1942 329
rect 1930 326 1938 328
rect 889 268 923 272
rect 1811 267 1874 275
rect 1847 246 1864 249
rect 905 241 916 245
rect 913 69 916 241
rect 1839 198 1850 201
rect 1856 160 1860 165
rect 1826 156 1860 160
rect 913 65 915 69
rect 1858 61 1864 64
rect 890 43 931 50
rect 913 8 916 38
rect 913 5 1094 8
rect 1091 1 1094 5
rect 1091 -2 1799 1
rect 1796 -3 1915 -2
rect 1923 -3 1924 -2
rect 1796 -5 1924 -3
rect 1911 -6 1926 -5
rect 1899 -12 1902 -8
rect 1735 -15 1906 -12
<< metal2 >>
rect 1820 326 1926 329
rect 1820 241 1823 326
rect 1813 198 1835 201
rect 905 156 911 159
rect 898 -4 901 82
rect 908 4 911 156
rect 1843 81 1846 246
rect 1854 198 1867 201
rect 1820 78 1846 81
rect 916 39 919 65
rect 1858 61 1864 64
rect 908 1 1090 4
rect 1087 -4 1090 1
rect 898 -7 1083 -4
rect 1087 -7 1789 -4
rect 1080 -12 1083 -7
rect 1080 -15 1731 -12
rect 1786 -19 1789 -7
rect 1857 -19 1860 61
rect 1786 -22 1860 -19
<< polycontact >>
rect 1938 324 1942 328
rect 1864 245 1868 249
rect 1856 165 1860 169
rect 1864 61 1868 65
rect 1924 -5 1928 -1
rect 1902 -12 1906 -8
<< m2contact >>
rect 1926 326 1930 330
rect 1843 246 1847 250
rect 901 156 905 160
rect 1809 198 1813 202
rect 1835 198 1839 202
rect 1850 198 1854 202
rect 915 65 919 69
rect 1854 61 1858 65
rect 916 35 920 39
rect 1731 -15 1735 -11
use totdiff3  totdiff3_0
timestamp 1523170410
transform 1 0 -507 0 1 672
box 507 -672 1412 -374
use totdiff3  totdiff3_1
timestamp 1523170410
transform 1 0 415 0 1 672
box 507 -672 1412 -374
use comp  comp_0
timestamp 1523170410
transform 1 0 1886 0 1 240
box -22 -240 296 83
<< end >>
