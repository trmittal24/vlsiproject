* Wed Feb 28 17:04:02 CET 2007
.subckt nd3v5x6 a b c vdd vss z
*SPICE circuit <nd3v5x6> from XCircuit v3.4 rev 26

m1 z c vdd vdd p w=81u l=2u ad='81u*5u+12p' as='81u*5u+12p' pd='81u*2+14u' ps='81u*2+14u'
m2 z a vdd vdd p w=81u l=2u ad='81u*5u+12p' as='81u*5u+12p' pd='81u*2+14u' ps='81u*2+14u'
m3 n1 a vss vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m4 n2 b n1 vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m5 z c n2 vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m6 z b vdd vdd p w=81u l=2u ad='81u*5u+12p' as='81u*5u+12p' pd='81u*2+14u' ps='81u*2+14u'
.ends
