* Spice description of an2_x2
* Spice driver version 134999461
* Date 31/05/2007 at 21:32:16
* vxlib 0.13um values
.subckt an2_x2 a b vdd vss z
M1a vdd   a     zn    vdd p  L=0.12U  W=1.375U AS=0.364375P AD=0.364375P PS=3.28U   PD=3.28U
M1b zn    b     vdd   vdd p  L=0.12U  W=1.375U AS=0.364375P AD=0.364375P PS=3.28U   PD=3.28U
M1z z     zn    vdd   vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M2a sig2  a     vss   vss n  L=0.12U  W=1.155U AS=0.306075P AD=0.306075P PS=2.84U   PD=2.84U
M2b zn    b     sig2  vss n  L=0.12U  W=1.155U AS=0.306075P AD=0.306075P PS=2.84U   PD=2.84U
M2z vss   zn    z     vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
C6  a     vss   0.543f
C7  b     vss   0.625f
C4  z     vss   0.790f
C1  zn    vss   0.766f
.ends
