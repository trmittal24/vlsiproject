* Spice description of xor2_x05
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:11
*
.subckt xor2_x05 a b vdd vss z 
M3  sig4  a     vdd   vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M4  vdd   b     sig5  vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M2  z     sig5  sig4  vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M1  sig5  sig4  z     vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M5  sig2  sig4  vss   vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M6  z     sig5  sig2  vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M7  sig4  b     z     vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M8  vss   a     sig4  vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M9  sig5  b     vss   vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
C8  a     vss   1.334f
C7  b     vss   1.249f
C6  vdd   vss   1.535f
C5  sig5  vss   2.265f
C4  sig4  vss   1.383f
C1  z     vss   2.558f
.ends
