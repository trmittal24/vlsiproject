* SPICE3 file created from counter.ext - technology: scmos

.include t14y_tsmc_025_level3.txt

.option scale=1u

M1000 t_0_cp an2v0x3_0_zn t_2_vdd t_2_vdd cmosp w=20 l=2
+ ad=160 pd=56 as=3514 ps=1266 
M1001 t_2_vdd an2v0x3_0_zn t_0_cp t_2_vdd cmosp w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1002 an2v0x3_0_zn an2v0x3_0_a t_2_vdd t_2_vdd cmosp w=20 l=2
+ ad=166 pd=62 as=0 ps=0 
M1003 t_2_vdd an2v0x3_0_b an2v0x3_0_zn t_2_vdd cmosp w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1004 t_2_vss an2v0x3_0_zn t_0_cp t_2_vss cmosn w=20 l=2
+ ad=2497 pd=1052 as=126 ps=54 
M1005 an2v0x3_0_a_30_9# an2v0x3_0_a t_2_vss t_2_vss cmosn w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1006 an2v0x3_0_zn an2v0x3_0_b an2v0x3_0_a_30_9# t_2_vss cmosn w=17 l=2
+ ad=97 pd=48 as=0 ps=0 
M1007 t_2_vdd t_0_d t_0_z t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=168 ps=70 
M1008 t_0_d t_0_n4 t_2_vdd t_2_vdd cmosp w=14 l=2
+ ad=82 pd=42 as=0 ps=0 
M1009 t_0_a_44_52# t_0_d t_2_vdd t_2_vdd cmosp w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1010 t_0_n4 t_0_ci t_0_a_44_52# t_2_vdd cmosp w=6 l=2
+ ad=78 pd=40 as=0 ps=0 
M1011 t_0_n2 t_0_cn t_0_n4 t_2_vdd cmosp w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1012 t_2_vdd t_0_n1 t_0_n2 t_2_vdd cmosp w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1013 t_0_a_81_58# t_0_n2 t_2_vdd t_2_vdd cmosp w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1014 t_0_n1 t_0_cn t_0_a_81_58# t_2_vdd cmosp w=6 l=2
+ ad=83 pd=42 as=0 ps=0 
M1015 t_2_vss t_0_d t_0_z t_2_vss cmosn w=14 l=2
+ ad=0 pd=0 as=82 ps=42 
M1016 t_2_vss t_0_n4 t_0_d t_2_vss cmosn w=7 l=2
+ ad=0 pd=0 as=47 ps=28 
M1017 t_0_a_98_51# t_0_ci t_0_n1 t_2_vdd cmosp w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1018 t_2_vdd t_0_d t_0_a_98_51# t_2_vdd cmosp w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1019 t_0_ci t_0_cn t_2_vdd t_2_vdd cmosp w=11 l=2
+ ad=67 pd=36 as=0 ps=0 
M1020 t_0_cn t_0_cp t_2_vdd t_2_vdd cmosp w=10 l=2
+ ad=62 pd=34 as=0 ps=0 
M1021 t_2_vss t_0_cn t_0_ci t_2_vss cmosn w=6 l=2
+ ad=0 pd=0 as=42 ps=26 
M1022 t_0_a_44_17# t_0_d t_2_vss t_2_vss cmosn w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1023 t_0_n4 t_0_cn t_0_a_44_17# t_2_vss cmosn w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1024 t_0_n2 t_0_ci t_0_n4 t_2_vss cmosn w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1025 t_2_vss t_0_n1 t_0_n2 t_2_vss cmosn w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1026 t_0_a_81_17# t_0_n2 t_2_vss t_2_vss cmosn w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1027 t_0_n1 t_0_ci t_0_a_81_17# t_2_vss cmosn w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1028 t_0_a_98_17# t_0_cn t_0_n1 t_2_vss cmosn w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1029 t_2_vss t_0_d t_0_a_98_17# t_2_vss cmosn w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1030 t_0_cn t_0_cp t_2_vss t_2_vss cmosn w=7 l=2
+ ad=49 pd=28 as=0 ps=0 
M1031 xor2v0x3_0_bn xor2v0x3_1_b t_2_vdd t_2_vdd cmosp w=28 l=2
+ ad=672 pd=216 as=0 ps=0 
M1032 t_2_vdd xor2v0x3_1_b xor2v0x3_0_bn t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1033 xor2v0x3_0_bn xor2v0x3_1_b t_2_vdd t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1034 t_1_cp xor2v0x3_0_an xor2v0x3_0_bn t_2_vdd cmosp w=28 l=2
+ ad=582 pd=216 as=0 ps=0 
M1035 xor2v0x3_0_an xor2v0x3_0_bn t_1_cp t_2_vdd cmosp w=13 l=2
+ ad=494 pd=184 as=0 ps=0 
M1036 t_1_cp xor2v0x3_0_bn xor2v0x3_0_an t_2_vdd cmosp w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1037 xor2v0x3_0_bn xor2v0x3_0_an t_1_cp t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1038 t_1_cp xor2v0x3_0_an xor2v0x3_0_bn t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1039 xor2v0x3_0_an xor2v0x3_0_bn t_1_cp t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1040 t_2_vdd t_0_z xor2v0x3_0_an t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1041 xor2v0x3_0_an t_0_z t_2_vdd t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1042 xor2v0x3_0_bn xor2v0x3_1_b t_2_vss t_2_vss cmosn w=11 l=2
+ ad=118 pd=50 as=0 ps=0 
M1043 t_2_vss xor2v0x3_1_b xor2v0x3_0_bn t_2_vss cmosn w=17 l=2
+ ad=0 pd=0 as=0 ps=0 
M1044 xor2v0x3_0_an xor2v0x3_1_b t_1_cp t_2_vss cmosn w=14 l=2
+ ad=224 pd=88 as=342 ps=148 
M1045 t_1_cp xor2v0x3_1_b xor2v0x3_0_an t_2_vss cmosn w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1046 xor2v0x3_0_a_61_7# xor2v0x3_0_an t_1_cp t_2_vss cmosn w=19 l=2
+ ad=95 pd=48 as=0 ps=0 
M1047 t_2_vss xor2v0x3_0_bn xor2v0x3_0_a_61_7# t_2_vss cmosn w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1048 xor2v0x3_0_a_80_7# xor2v0x3_0_bn t_2_vss t_2_vss cmosn w=19 l=2
+ ad=95 pd=48 as=0 ps=0 
M1049 t_1_cp xor2v0x3_0_an xor2v0x3_0_a_80_7# t_2_vss cmosn w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1050 xor2v0x3_0_an t_0_z t_2_vss t_2_vss cmosn w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1051 t_2_vss t_0_z xor2v0x3_0_an t_2_vss cmosn w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1052 t_2_vdd t_1_d t_1_z t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=168 ps=70 
M1053 t_1_d t_1_n4 t_2_vdd t_2_vdd cmosp w=14 l=2
+ ad=82 pd=42 as=0 ps=0 
M1054 t_1_a_44_52# t_1_d t_2_vdd t_2_vdd cmosp w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1055 t_1_n4 t_1_ci t_1_a_44_52# t_2_vdd cmosp w=6 l=2
+ ad=78 pd=40 as=0 ps=0 
M1056 t_1_n2 t_1_cn t_1_n4 t_2_vdd cmosp w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1057 t_2_vdd t_1_n1 t_1_n2 t_2_vdd cmosp w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1058 t_1_a_81_58# t_1_n2 t_2_vdd t_2_vdd cmosp w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1059 t_1_n1 t_1_cn t_1_a_81_58# t_2_vdd cmosp w=6 l=2
+ ad=83 pd=42 as=0 ps=0 
M1060 t_2_vss t_1_d t_1_z t_2_vss cmosn w=14 l=2
+ ad=0 pd=0 as=82 ps=42 
M1061 t_2_vss t_1_n4 t_1_d t_2_vss cmosn w=7 l=2
+ ad=0 pd=0 as=47 ps=28 
M1062 t_1_a_98_51# t_1_ci t_1_n1 t_2_vdd cmosp w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1063 t_2_vdd t_1_d t_1_a_98_51# t_2_vdd cmosp w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1064 t_1_ci t_1_cn t_2_vdd t_2_vdd cmosp w=11 l=2
+ ad=67 pd=36 as=0 ps=0 
M1065 t_1_cn t_1_cp t_2_vdd t_2_vdd cmosp w=10 l=2
+ ad=62 pd=34 as=0 ps=0 
M1066 t_2_vss t_1_cn t_1_ci t_2_vss cmosn w=6 l=2
+ ad=0 pd=0 as=42 ps=26 
M1067 t_1_a_44_17# t_1_d t_2_vss t_2_vss cmosn w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1068 t_1_n4 t_1_cn t_1_a_44_17# t_2_vss cmosn w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1069 t_1_n2 t_1_ci t_1_n4 t_2_vss cmosn w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1070 t_2_vss t_1_n1 t_1_n2 t_2_vss cmosn w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1071 t_1_a_81_17# t_1_n2 t_2_vss t_2_vss cmosn w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1072 t_1_n1 t_1_ci t_1_a_81_17# t_2_vss cmosn w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1073 t_1_a_98_17# t_1_cn t_1_n1 t_2_vss cmosn w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1074 t_2_vss t_1_d t_1_a_98_17# t_2_vss cmosn w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1075 t_1_cn t_1_cp t_2_vss t_2_vss cmosn w=7 l=2
+ ad=49 pd=28 as=0 ps=0 
M1076 xor2v0x3_1_bn xor2v0x3_1_b t_2_vdd t_2_vdd cmosp w=28 l=2
+ ad=672 pd=216 as=0 ps=0 
M1077 t_2_vdd xor2v0x3_1_b xor2v0x3_1_bn t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1078 xor2v0x3_1_bn xor2v0x3_1_b t_2_vdd t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1079 t_2_cp xor2v0x3_1_an xor2v0x3_1_bn t_2_vdd cmosp w=28 l=2
+ ad=582 pd=216 as=0 ps=0 
M1080 xor2v0x3_1_an xor2v0x3_1_bn t_2_cp t_2_vdd cmosp w=13 l=2
+ ad=494 pd=184 as=0 ps=0 
M1081 t_2_cp xor2v0x3_1_bn xor2v0x3_1_an t_2_vdd cmosp w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1082 xor2v0x3_1_bn xor2v0x3_1_an t_2_cp t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1083 t_2_cp xor2v0x3_1_an xor2v0x3_1_bn t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1084 xor2v0x3_1_an xor2v0x3_1_bn t_2_cp t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1085 t_2_vdd t_1_z xor2v0x3_1_an t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1086 xor2v0x3_1_an t_1_z t_2_vdd t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1087 xor2v0x3_1_bn xor2v0x3_1_b t_2_vss t_2_vss cmosn w=11 l=2
+ ad=118 pd=50 as=0 ps=0 
M1088 t_2_vss xor2v0x3_1_b xor2v0x3_1_bn t_2_vss cmosn w=17 l=2
+ ad=0 pd=0 as=0 ps=0 
M1089 xor2v0x3_1_an xor2v0x3_1_b t_2_cp t_2_vss cmosn w=14 l=2
+ ad=224 pd=88 as=342 ps=148 
M1090 t_2_cp xor2v0x3_1_b xor2v0x3_1_an t_2_vss cmosn w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1091 xor2v0x3_1_a_61_7# xor2v0x3_1_an t_2_cp t_2_vss cmosn w=19 l=2
+ ad=95 pd=48 as=0 ps=0 
M1092 t_2_vss xor2v0x3_1_bn xor2v0x3_1_a_61_7# t_2_vss cmosn w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1093 xor2v0x3_1_a_80_7# xor2v0x3_1_bn t_2_vss t_2_vss cmosn w=19 l=2
+ ad=95 pd=48 as=0 ps=0 
M1094 t_2_cp xor2v0x3_1_an xor2v0x3_1_a_80_7# t_2_vss cmosn w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1095 xor2v0x3_1_an t_1_z t_2_vss t_2_vss cmosn w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1096 t_2_vss t_1_z xor2v0x3_1_an t_2_vss cmosn w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1097 t_2_vdd t_2_d t_2_z t_2_vdd cmosp w=28 l=2
+ ad=0 pd=0 as=168 ps=70 
M1098 t_2_d t_2_n4 t_2_vdd t_2_vdd cmosp w=14 l=2
+ ad=82 pd=42 as=0 ps=0 
M1099 t_2_a_44_52# t_2_d t_2_vdd t_2_vdd cmosp w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1100 t_2_n4 t_2_ci t_2_a_44_52# t_2_vdd cmosp w=6 l=2
+ ad=78 pd=40 as=0 ps=0 
M1101 t_2_n2 t_2_cn t_2_n4 t_2_vdd cmosp w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1102 t_2_vdd t_2_n1 t_2_n2 t_2_vdd cmosp w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1103 t_2_a_81_58# t_2_n2 t_2_vdd t_2_vdd cmosp w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1104 t_2_n1 t_2_cn t_2_a_81_58# t_2_vdd cmosp w=6 l=2
+ ad=83 pd=42 as=0 ps=0 
M1105 t_2_vss t_2_d t_2_z t_2_vss cmosn w=14 l=2
+ ad=0 pd=0 as=82 ps=42 
M1106 t_2_vss t_2_n4 t_2_d t_2_vss cmosn w=7 l=2
+ ad=0 pd=0 as=47 ps=28 
M1107 t_2_a_98_51# t_2_ci t_2_n1 t_2_vdd cmosp w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1108 t_2_vdd t_2_d t_2_a_98_51# t_2_vdd cmosp w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1109 t_2_ci t_2_cn t_2_vdd t_2_vdd cmosp w=11 l=2
+ ad=67 pd=36 as=0 ps=0 
M1110 t_2_cn t_2_cp t_2_vdd t_2_vdd cmosp w=10 l=2
+ ad=62 pd=34 as=0 ps=0 
M1111 t_2_vss t_2_cn t_2_ci t_2_vss cmosn w=6 l=2
+ ad=0 pd=0 as=42 ps=26 
M1112 t_2_a_44_17# t_2_d t_2_vss t_2_vss cmosn w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1113 t_2_n4 t_2_cn t_2_a_44_17# t_2_vss cmosn w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1114 t_2_n2 t_2_ci t_2_n4 t_2_vss cmosn w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1115 t_2_vss t_2_n1 t_2_n2 t_2_vss cmosn w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1116 t_2_a_81_17# t_2_n2 t_2_vss t_2_vss cmosn w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1117 t_2_n1 t_2_ci t_2_a_81_17# t_2_vss cmosn w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1118 t_2_a_98_17# t_2_cn t_2_n1 t_2_vss cmosn w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1119 t_2_vss t_2_d t_2_a_98_17# t_2_vss cmosn w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1120 t_2_cn t_2_cp t_2_vss t_2_vss cmosn w=7 l=2
+ ad=49 pd=28 as=0 ps=0 
C0 t_2_vss t_0_cn 17.1fF
C1 t_2_vdd t_1_z 11.0fF
C2 t_2_n4 t_2_vss 7.3fF
C3 t_0_d t_2_vss 28.2fF
C4 t_1_n2 t_2_vdd 12.4fF
C5 t_2_vss t_1_d 28.2fF
C6 t_2_ci t_2_vss 27.5fF
C7 t_1_ci t_1_d 4.2fF
C8 t_2_vdd t_0_cn 46.5fF
C9 t_2_n4 t_2_vdd 8.9fF
C10 t_1_cn t_2_vss 17.1fF
C11 t_0_d t_2_vdd 18.0fF
C12 t_0_ci t_2_vss 27.5fF
C13 t_2_cp t_2_vss 9.0fF
C14 t_1_d t_2_vdd 18.0fF
C15 t_2_ci t_2_vdd 16.6fF
C16 t_2_vss t_1_n4 7.3fF
C17 t_2_cn t_2_vss 17.1fF
C18 xor2v0x3_0_an t_2_vss 18.3fF
C19 t_1_cn t_2_vdd 46.5fF
C20 t_0_ci t_2_vdd 16.6fF
C21 t_2_n2 t_2_vss 7.2fF
C22 t_1_ci t_2_vss 27.5fF
C23 t_2_cp t_2_vdd 23.0fF
C24 t_2_ci t_2_d 4.2fF
C25 t_1_n4 t_2_vdd 8.9fF
C26 t_2_cn t_2_vdd 46.5fF
C27 xor2v0x3_0_an t_2_vdd 19.1fF
C28 t_2_vss xor2v0x3_0_bn 12.6fF
C29 t_2_n2 t_2_vdd 12.4fF
C30 t_0_z t_2_vss 12.2fF
C31 t_1_ci t_2_vdd 16.6fF
C32 t_2_vss an2v0x3_0_zn 9.5fF
C33 xor2v0x3_1_an t_2_cp 3.6fF
C34 t_2_cp xor2v0x3_1_b 6.8fF
C35 xor2v0x3_0_bn t_2_vdd 24.1fF
C36 t_2_vss t_2_d 28.2fF
C37 t_2_n1 t_2_vss 9.9fF
C38 xor2v0x3_1_an t_2_vss 18.3fF
C39 t_0_z t_2_vdd 11.0fF
C40 t_2_vss xor2v0x3_1_b 51.1fF
C41 an2v0x3_0_zn t_2_vdd 13.3fF
C42 t_2_vss t_0_n4 7.3fF
C43 t_2_d t_2_vdd 18.0fF
C44 t_2_n1 t_2_vdd 8.4fF
C45 an2v0x3_0_b t_2_vss 5.5fF
C46 t_2_z t_2_vdd 2.7fF
C47 t_1_n1 t_2_vss 9.9fF
C48 xor2v0x3_1_an t_2_vdd 19.1fF
C49 xor2v0x3_1_b t_2_vdd 38.6fF
C50 t_0_n4 t_2_vdd 8.9fF
C51 t_2_vss an2v0x3_0_a 6.3fF
C52 an2v0x3_0_b t_2_vdd 6.5fF
C53 t_1_n1 t_2_vdd 8.4fF
C54 xor2v0x3_0_an t_1_cp 3.6fF
C55 t_1_cp t_2_vss 9.0fF
C56 t_2_vss t_0_cp 4.7fF
C57 an2v0x3_0_a t_2_vdd 5.3fF
C58 xor2v0x3_1_bn t_2_cp 8.8fF
C59 t_1_cp xor2v0x3_0_bn 7.1fF
C60 t_1_cp t_2_vdd 22.3fF
C61 t_0_cp t_2_vdd 18.8fF
C62 xor2v0x3_1_bn t_2_vss 12.6fF
C63 t_2_vss t_0_n1 9.9fF
C64 t_2_vss t_0_n2 7.2fF
C65 t_2_vss t_1_z 12.1fF
C66 t_0_d t_0_ci 4.2fF
C67 xor2v0x3_1_bn t_2_vdd 24.1fF
C68 t_0_n1 t_2_vdd 8.4fF
C69 t_2_vss t_1_n2 7.2fF
C70 t_0_n2 t_2_vdd 12.4fF
C71 t_2_vss 0 7.5fF
C72 t_2_vdd 0 7.9fF


v_dd t_2_vdd 0 5
v_ss t_2_vss 0 0
v_gg_cp an2v0x3_0_a 0 PULSE(0 5 0 0.1n 0.1n 15n 30n)
*v_gg_t b 0 PULSE(5 0 10n 0 0 20n 500n)
v_dd_en an2v0x3_0_b 0 5
v_dd_ud xor2v0x3_1_b 0 5

.control
 tran 0.01n 300n
 plot (an2v0x3_0_a + 5) (t_0_z) (t_1_z - 5) (t_2_z - 10)
.endc

.end