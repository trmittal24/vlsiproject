* Spice description of cgi2_x05
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:09
*
.subckt cgi2_x05 a b c vdd vss z 
M04 n2    b     vdd   vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M05 z     c     n2    vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M01 vdd   a     sig5  vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M03 sig5  b     z     vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M02 n2    a     vdd   vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M07 vss   a     sig2  vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M06 n3    a     vss   vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M08 z     b     n3    vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M09 vss   b     sig2  vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M10 sig2  c     z     vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
C10 c     vss   1.014f
C9  b     vss   2.187f
C8  a     vss   1.308f
C7  vdd   vss   1.521f
C6  n2    vss   0.807f
C4  z     vss   1.920f
C2  sig2  vss   1.085f
.ends
