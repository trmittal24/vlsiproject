magic
tech scmos
timestamp 1523178222
<< error_s >>
rect 1886 -182 1887 -181
<< polysilicon >>
rect 1939 313 1941 324
rect 1868 246 1901 248
rect 1860 166 1903 168
rect 1967 85 1969 89
rect 1897 83 1969 85
rect 1897 64 1899 83
rect 1868 62 1899 64
rect 1903 -8 1905 9
rect 1925 -1 1927 8
rect 1925 -6 1927 -5
<< metal1 >>
rect 1930 328 1942 329
rect 1930 326 1938 328
rect 1811 267 1874 275
rect 1847 246 1864 249
rect 1819 189 1823 245
rect 1839 198 1850 201
rect 1856 160 1860 165
rect 1826 156 1856 160
rect 922 -45 925 118
rect 1823 93 1838 97
rect 1835 74 1838 93
rect 1826 70 1838 74
rect 1809 44 1820 51
rect 1817 -57 1820 44
rect 1826 43 1830 70
rect 2179 68 2189 75
rect 1842 61 1864 64
rect 1826 39 1863 43
rect 1813 -61 1820 -57
rect 1824 -3 1915 -2
rect 1923 -3 1924 -2
rect 1824 -5 1924 -3
rect 1813 -106 1816 -61
rect 1824 -76 1827 -5
rect 1911 -6 1926 -5
rect 1831 -11 1902 -8
rect 1831 -82 1834 -11
rect 1920 -19 1923 -6
rect 1897 -22 1923 -19
rect 1897 -36 1900 -22
rect 1961 -32 1970 9
rect 2185 -11 2189 68
rect 2186 -36 2189 -11
rect 1988 -39 2190 -36
rect 1810 -114 1816 -106
rect 1809 -118 1816 -114
rect 1824 -85 1834 -82
rect 1985 -43 2190 -39
rect 1824 -125 1827 -85
rect 1985 -104 1989 -43
rect 1980 -111 1989 -104
rect 1980 -112 1988 -111
rect 1824 -128 1836 -125
rect 1833 -235 1836 -128
rect 1866 -181 1887 -177
rect 1871 -182 1884 -181
rect 1883 -235 1887 -185
rect 1825 -239 1887 -235
<< metal2 >>
rect 1820 326 1926 329
rect 1820 241 1823 326
rect 1813 198 1835 201
rect 1819 97 1823 185
rect 1843 81 1846 246
rect 1854 198 1867 201
rect 1820 78 1849 81
rect 1838 -82 1841 61
rect 1824 -85 1841 -82
rect 1824 -157 1827 -85
rect 1846 -93 1849 78
rect 1856 -83 1859 156
rect 1863 -73 1866 39
rect 1872 -73 1885 -72
rect 1863 -76 1891 -73
rect 1856 -87 1891 -83
rect 1885 -92 1891 -91
rect 1885 -93 1892 -92
rect 1846 -94 1892 -93
rect 1846 -96 1895 -94
rect 1871 -97 1884 -96
rect 1827 -161 1847 -157
rect 1843 -177 1847 -161
rect 1843 -181 1862 -177
<< polycontact >>
rect 1938 324 1942 328
rect 1864 245 1868 249
rect 1856 165 1860 169
rect 1864 61 1868 65
rect 1924 -5 1928 -1
rect 1902 -12 1906 -8
<< m2contact >>
rect 1926 326 1930 330
rect 1843 246 1847 250
rect 1809 198 1813 202
rect 1835 198 1839 202
rect 1850 198 1854 202
rect 1819 185 1823 189
rect 1856 156 1860 160
rect 1819 93 1823 97
rect 1838 61 1842 65
rect 1863 39 1867 43
rect 1823 -161 1827 -157
rect 1862 -181 1866 -177
use totdiff3  totdiff3_1
timestamp 1523176862
transform 1 0 415 0 1 672
box 507 -672 1412 -374
use comp  comp_0
timestamp 1523176862
transform 1 0 1886 0 1 240
box -22 -240 296 83
use totdiff3  totdiff3_0
timestamp 1523176862
transform 1 0 415 0 1 355
box 507 -672 1412 -374
use mux  mux_0
timestamp 1523176862
transform 1 0 1915 0 1 -103
box -29 -160 85 80
<< end >>
