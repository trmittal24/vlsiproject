* Spice description of oai22_x2
* Spice driver version 134999461
* Date 31/05/2007 at 21:35:23
* vxlib 0.13um values
.subckt oai22_x2 a1 a2 b1 b2 vdd vss z
M1a vdd   a1    sig6  vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M1b n1b   a1    vdd   vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M2a sig6  a2    z     vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M2b z     a2    n1b   vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M3a vdd   b1    n2a   vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M3b n2b   b1    vdd   vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M4a n2a   b2    z     vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M4b z     b2    n2b   vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M5  vss   a1    sig2  vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M6  sig2  a2    vss   vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M7  sig2  b1    z     vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M8  z     b2    sig2  vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
C9  a1    vss   0.915f
C12 a2    vss   0.584f
C10 b1    vss   0.966f
C8  b2    vss   0.659f
C2  sig2  vss   0.451f
C3  z     vss   1.810f
.ends
