* Mon Apr 30 10:20:21 CEST 2007
.subckt xor2v8x05 a b vdd vss z
*SPICE circuit <xor2v8x05> from XCircuit v3.4 rev 26

m1 z zn vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m2 z zn vdd vdd p w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m3 an b zn vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m4 zn bn an vdd p w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m5 bn b vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m6 bn b vdd vdd p w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m7 an a vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m8 ai an vdd vdd p w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m9 ai an vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m10 ai bn zn vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m11 an a vdd vdd p w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m12 zn b ai vdd p w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
.ends
