* Tue Dec 14 18:00:47 CET 2004
.subckt xoon21v0x1 a1 a2 b vdd vss z 
*SPICE circuit <xoon21v0x1> from XCircuit v3.20

m1 an a1 vss vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m2 an a2 vss vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m3 n1 a1 vdd vdd p w=49u l=2.3636u ad='49u*5u+12p' as='49u*5u+12p' pd='49u*2+14u' ps='49u*2+14u'
m4 an a2 n1 vdd p w=49u l=2.3636u ad='49u*5u+12p' as='49u*5u+12p' pd='49u*2+14u' ps='49u*2+14u'
m5 z bn an vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m6 bn b vss vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m7 n2 an vss vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m8 z bn n2 vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m9 bn b vdd vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m10 z b an vss n w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m11 z an bn vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
.ends
