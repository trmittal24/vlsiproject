* Spice description of aoi21_x05
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:09
*
.subckt aoi21_x05 a1 a2 b vdd vss z 
M3  z     b     sig4  vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M2  sig4  a2    vdd   vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M1  vdd   a1    sig4  vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M6  z     b     vss   vss n  L=0.13U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U  
M5  sig3  a2    z     vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M4  vss   a1    sig3  vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
C8  a1    vss   1.046f
C7  b     vss   1.632f
C6  a2    vss   1.035f
C5  vdd   vss   1.114f
C4  sig4  vss   0.529f
C1  z     vss   2.253f
.ends
