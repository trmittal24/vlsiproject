* Thu Jan 27 22:08:39 CET 2005
.subckt nr2v0x3 a b vdd vss z 
*SPICE circuit <nr2v0x3> from XCircuit v3.10

m1 z a vss vss n w=23u l=2.3636u ad='23u*5u+12p' as='23u*5u+12p' pd='23u*2+14u' ps='23u*2+14u'
m2 n1 a vdd vdd p w=84u l=2.3636u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m3 z b vss vss n w=23u l=2.3636u ad='23u*5u+12p' as='23u*5u+12p' pd='23u*2+14u' ps='23u*2+14u'
m4 z b n1 vdd p w=84u l=2.3636u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
.ends
