* Sat Apr  9 11:13:33 CEST 2005
.subckt nr2av0x6 a b vdd vss z 
*SPICE circuit <nr2av0x6> from XCircuit v3.20

m1 an a vss vss n w=24u l=2u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m2 an a vdd vdd p w=48u l=2u ad='48u*5u+12p' as='48u*5u+12p' pd='48u*2+14u' ps='48u*2+14u'
m3 z an vss vss n w=45u l=2u ad='45u*5u+12p' as='45u*5u+12p' pd='45u*2+14u' ps='45u*2+14u'
m4 n1 an vdd vdd p w=168u l=2u ad='168u*5u+12p' as='168u*5u+12p' pd='168u*2+14u' ps='168u*2+14u'
m5 z b vss vss n w=45u l=2u ad='45u*5u+12p' as='45u*5u+12p' pd='45u*2+14u' ps='45u*2+14u'
m6 z b n1 vdd p w=168u l=2u ad='168u*5u+12p' as='168u*5u+12p' pd='168u*2+14u' ps='168u*2+14u'
.ends
