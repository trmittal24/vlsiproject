* Spice description of vfeed1
* Spice driver version 134999461
* Date 31/05/2007 at 21:35:53
* vxlib 0.13um values
.subckt vfeed1 vdd vss
.ends
