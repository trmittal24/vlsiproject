* Mon Aug 16 14:10:57 CEST 2004
.subckt aoi31v0x1 a1 a2 a3 b vdd vss z 
*SPICE circuit <aoi31v0x1> from XCircuit v3.10

m1 n1 a1 vss vss n w=17u l=2.3636u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m2 n3 a1 vdd vdd p w=27u l=2.3636u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
m3 n3 a3 vdd vdd p w=27u l=2.3636u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
m4 n3 a2 vdd vdd p w=27u l=2.3636u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
m5 n2 a2 n1 vss n w=17u l=2.3636u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m6 z b vss vss n w=7u l=2.3636u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m7 z a3 n2 vss n w=17u l=2.3636u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m8 z b n3 vdd p w=27u l=2.3636u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
.ends
