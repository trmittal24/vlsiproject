* Spice description of vsstie
* Spice driver version 134999461
* Date  6/02/2007 at 12:04:04
* rgalib 0.13um values
.subckt vsstie vdd vss z
Mtr_00001 z     vdd   vss   vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00002 vss   vdd   z     vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00003 z     vdd   sig5  vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
Mtr_00004 sig4  vdd   z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
C1  z     vss   0.660f
.ends
