* Spice description of aoi22_x2
* Spice driver version 134999461
* Date 22/07/2007 at 10:57:25
* vsxlib 0.13um values
.subckt aoi22_x2 a1 a2 b1 b2 vdd vss z
M1a vdd   a1    4a    vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M1b 4a    a1    vdd   vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M2a 4a    a2    vdd   vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M2b vdd   a2    4a    vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M3a z     b1    4a    vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M3b 4a    b1    z     vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M4a 4a    b2    z     vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M4b z     b2    4a    vdd p  L=0.12U  W=2.035U AS=0.539275P AD=0.539275P PS=4.6U    PD=4.6U
M5  vss   a1    n1    vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M6  n1    a2    z     vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M7  n2    b1    vss   vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M8  z     b2    n2    vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
C9  4a    vss   0.956f
C8  a1    vss   0.662f
C6  a2    vss   0.942f
C5  b1    vss   0.644f
C4  b2    vss   0.910f
C1  z     vss   1.802f
.ends
