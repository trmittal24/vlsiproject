* Spice description of o4_x2
* Spice driver version 134999461
* Date 31/05/2007 at 10:39:38
* ssxlib 0.13um values
.subckt o4_x2 i0 i1 i2 i3 q vdd vss
Mtr_00001 sig2  i2    vss   vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
Mtr_00002 vss   i3    sig2  vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00003 vss   i0    sig2  vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00004 sig2  i1    vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00005 q     sig2  vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00006 sig8  i3    sig2  vdd p  L=0.12U  W=1.595U AS=0.422675P AD=0.422675P PS=3.72U   PD=3.72U
Mtr_00007 sig9  i1    sig8  vdd p  L=0.12U  W=1.595U AS=0.422675P AD=0.422675P PS=3.72U   PD=3.72U
Mtr_00008 sig11 i0    sig9  vdd p  L=0.12U  W=1.595U AS=0.422675P AD=0.422675P PS=3.72U   PD=3.72U
Mtr_00009 vdd   i2    sig11 vdd p  L=0.12U  W=1.595U AS=0.422675P AD=0.422675P PS=3.72U   PD=3.72U
Mtr_00010 vdd   sig2  q     vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
C7  i0    vss   0.684f
C4  i1    vss   0.646f
C6  i2    vss   0.683f
C3  i3    vss   0.624f
C5  q     vss   0.964f
C2  sig2  vss   1.098f
.ends
