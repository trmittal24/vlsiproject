* Spice description of aon21_x2
* Spice driver version 134999461
* Date 22/07/2007 at 10:57:29
* vsxlib 0.13um values
.subckt aon21_x2 a1 a2 b vdd vss z
M1  vdd   a1    3     vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M2  3     a2    vdd   vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M3_1 sig3  b     3     vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M3  z     sig3  vdd   vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M4  vss   a1    n1    vss n  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
M5_2 vss   sig3  z     vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
M5  n1    a2    sig3  vss n  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
M6  sig3  b     vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
C9  3     vss   0.198f
C7  a1    vss   0.647f
C6  a2    vss   0.568f
C5  b     vss   0.653f
C3  sig3  vss   0.638f
C2  z     vss   0.834f
.ends
