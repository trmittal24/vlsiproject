* Spice description of mxi2v2x05
* Spice driver version 134999461
* Date 17/05/2007 at  9:14:57
* wsclib 0.13um values
.subckt mxi2v2x05 a0 a1 s vdd vss z
M01 a0n   a0    vdd   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M02 a0n   a0    vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M03 vdd   a1    sig6  vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M04 vss   a1    sig6  vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M05 10    s     vdd   vdd p  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M06 10    s     vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M07 z     s     a0n   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M08 sig6  s     z     vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M09 sig6  10    z     vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M10 z     10    a0n   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
C5  10    vss   0.642f
C4  a0    vss   0.515f
C2  a0n   vss   0.255f
C7  a1    vss   0.408f
C8  s     vss   0.850f
C6  sig6  vss   0.244f
C3  z     vss   0.503f
.ends
