* Sat Aug 27 22:10:23 CEST 2005
.subckt iv1v5x3 a vdd vss z 
*SPICE circuit <iv1v5x3> from XCircuit v3.20

m1 z a vss vss n w=15u l=2.3636u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m2 z a vdd vdd p w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
.ends
