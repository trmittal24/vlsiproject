* functionality check of nd2av0x6, 0.13um, Berkeley generic bsim3 params
* nd2av0x6_func.cir 2007-08-29:12h15 graham
*
.include ../../../magic/subckt/vsclib013/spice_model.lib
.include ../../../magic/subckt/vsclib013/nd2av0x6.spi
.include ../../../magic/subckt/vsclib013/params.inc
*
x01 va   vb   vdd vss x01z nd2av0x6
x02 va   vb   vdd vss x02z nd2av0x6
*
.param unitcap=1.0f
cx01z  x01z  0 '6*unitcap'
cx02z  x02z  0 '130*6*unitcap'
* 
vdd vdd 0 'vdd'
vss 0 vss 'vss'
vstrobe strobe 0 dc 0 pulse (0 1 '0.97*tPER' '0.01*tPER' '0.01*tPER' '0.01*tPER' 'tPER')
*
* ba      00   10     11     01     00     01     11     10     00
*          0    1      0      1      0      1      0      1      0
*             thh_AZ thl_BZ tlh_AZ tll_BZ thh_BZ thl_AZ tlh_BZ tll_AZ
*                 0      1      2      3      4      5      6      7      8
Vb  vb 0 dc 0 pwl(0 'vss' '1*tPER' 'vss' '1*tPER+tRISE' 'vdd' '3*tPER' 'vdd' '3*tPER+tFALL' 'vss'
+           '4*tPER' 'vss' '4*tPER+tRISE' 'vdd' '6*tPER' 'vdd' '6*tPER+tFALL' 'vss' )
Va  va 0 dc 0 pwl(0 'vss' 'tRISE'  'vdd' '2*tPER' 'vdd'  '2*tPER+tFALL' 'vss'
+           '5*tPER' 'vss' '5*tPER+tRISE' 'vdd' '7*tPER' 'vdd' '7*tPER+tFALL' 'vss' )

.control
  set width=120 height=500 numdgt=3 noprintscale nobreak noaskquit=1
  tran $tstep 40000p
  linearize
  let a = va / $vdd
  let b = vb / $vdd
  let pa = va + ( $vdd + 0.3 )
  let pb = vb + 2 * ( $vdd + 0.3 )
  let pz = $vdd * (a or not (b)) - $vdd - 0.3
* check output is within 10mV of ideal at strobe point
  let perr =  vecmax ( pos ( abs (( pz - x02z + $vdd + 0.3 ) * strobe ) - 0.01 ))
  plot v(pa) v(pb) v(pz) v(x01z) v(x02z)
*  print col v(va) v(vb) v(x01z) v(x02z) > nd2av0x6_func.spo
  if perr > 0
    echo #Error: Functional simulation nd2av0x6_func.cir failed
    echo #Error: Functional simulation nd2av0x6_func.cir failed >> nd2av0x6_func.error
  else
    echo Functional simulation OK
  end
  destroy all
.endc
.end
