* Wed Apr  5 08:58:27 CEST 2006
.subckt bf1v0x6 a vdd vss z 
*SPICE circuit <bf1v0x6> from XCircuit v3.20

m1 an a vss vss n w=19u l=2u ad='19u*5u+12p' as='19u*5u+12p' pd='19u*2+14u' ps='19u*2+14u'
m2 an a vdd vdd p w=36u l=2u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
m3 z an vss vss n w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m4 z an vdd vdd p w=81u l=2u ad='81u*5u+12p' as='81u*5u+12p' pd='81u*2+14u' ps='81u*2+14u'
.ends
