* Spice description of on12_x4
* Spice driver version 134999461
* Date 21/07/2007 at 19:32:19
* sxlib 0.13um values
.subckt on12_x4 i0 i1 q vdd vss
Mtr_00001 vss   i0    sig3  vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00002 q     sig1  vss   vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00003 vss   sig1  q     vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00004 vss   sig3  sig1  vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00005 sig1  i1    vss   vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00006 vdd   i0    sig3  vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00007 sig6  sig3  sig1  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00008 vdd   sig1  q     vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00009 q     sig1  vdd   vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00010 vdd   i1    sig6  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
C8  i0    vss   1.016f
C7  i1    vss   0.908f
C4  q     vss   0.883f
C1  sig1  vss   0.928f
C3  sig3  vss   0.694f
.ends
