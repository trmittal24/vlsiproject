* Sat Aug 27 19:34:29 CEST 2005
.subckt nd2v4x3 a b vdd vss z 
*SPICE circuit <nd2v4x3> from XCircuit v3.20

m1 n1 a vss vss n w=19u l=2.3636u ad='19u*5u+12p' as='19u*5u+12p' pd='19u*2+14u' ps='19u*2+14u'
m2 z a vdd vdd p w=46u l=2.3636u ad='46u*5u+12p' as='46u*5u+12p' pd='46u*2+14u' ps='46u*2+14u'
m3 z b n1 vss n w=19u l=2.3636u ad='19u*5u+12p' as='19u*5u+12p' pd='19u*2+14u' ps='19u*2+14u'
m4 z b vdd vdd p w=46u l=2.3636u ad='46u*5u+12p' as='46u*5u+12p' pd='46u*2+14u' ps='46u*2+14u'
.ends
