* Wed Aug 31 12:58:40 CEST 2005
.subckt nd3v0x4 a b c vdd vss z 
*SPICE circuit <nd3v0x4> from XCircuit v3.20

m1 z c vdd vdd p w=50u l=2.3636u ad='50u*5u+12p' as='50u*5u+12p' pd='50u*2+14u' ps='50u*2+14u'
m2 z a vdd vdd p w=50u l=2.3636u ad='50u*5u+12p' as='50u*5u+12p' pd='50u*2+14u' ps='50u*2+14u'
m3 n1 a vss vss n w=50u l=2.3636u ad='50u*5u+12p' as='50u*5u+12p' pd='50u*2+14u' ps='50u*2+14u'
m4 n2 b n1 vss n w=50u l=2.3636u ad='50u*5u+12p' as='50u*5u+12p' pd='50u*2+14u' ps='50u*2+14u'
m5 z c n2 vss n w=50u l=2.3636u ad='50u*5u+12p' as='50u*5u+12p' pd='50u*2+14u' ps='50u*2+14u'
m6 z b vdd vdd p w=50u l=2.3636u ad='50u*5u+12p' as='50u*5u+12p' pd='50u*2+14u' ps='50u*2+14u'
.ends
