* Tue Aug 10 11:21:07 CEST 2004
.subckt nr2_x1 a b vdd vss z 
*SPICE circuit <nr2_x1> from XCircuit v3.10

m1 z a vss vss n w=11u l=2.3636u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m2 n1 a vdd vdd p w=39u l=2.3636u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m3 z b vss vss n w=11u l=2.3636u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m4 z b n1 vdd p w=39u l=2.3636u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
.ends
