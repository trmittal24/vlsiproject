* Tue Feb 20 08:57:11 CET 2007
.subckt iv1v0x2 a vdd vss z
*SPICE circuit <iv1v0x2> from XCircuit v3.4 rev 26

m1 z a vss vss n w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m2 z a vdd vdd p w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
.ends
