* Spice description of vsstie
* Spice driver version 134999461
* Date 17/06/2007 at 14:03:45
* vgalib 0.13um values
.subckt vsstie vdd vss z
Mtr_00001 z     sig3  vss   vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00002 vss   sig3  z     vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00003 vdd   z     sig3  vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
Mtr_00004 sig3  z     vdd   vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
C3  sig3  vss   0.732f
C1  z     vss   1.095f
.ends
