* Tue Feb 20 08:57:11 CET 2007
.subckt iv1v0x4 a vdd vss z
*SPICE circuit <iv1v0x4> from XCircuit v3.4 rev 26

m1 z a vss vss n w=36u l=2u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
m2 z a vdd vdd p w=52u l=2u ad='52u*5u+12p' as='52u*5u+12p' pd='52u*2+14u' ps='52u*2+14u'
.ends
