* Spice description of nr2av0x1
* Spice driver version 134999461
* Date 17/06/2007 at 14:03:20
* vgalib 0.13um values
.subckt nr2av0x1 a b vdd vss z
Mtr_00001 z     sig2  vss   vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00002 vss   b     z     vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00003 vss   vss   sig3  vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00004 sig2  a     vss   vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00005 z     b     sig9  vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
Mtr_00006 sig9  sig2  vdd   vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
Mtr_00007 sig2  a     vdd   vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
Mtr_00008 vdd   vdd   sig8  vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
C4  a     vss   0.508f
C6  b     vss   0.535f
C2  sig2  vss   0.815f
C5  z     vss   0.921f
.ends
