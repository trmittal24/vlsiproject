* Tue Dec 14 08:05:47 CET 2004
.subckt aoi211v0x2 a1 a2 b c vdd vss z 
*SPICE circuit <aoi211v0x2> from XCircuit v3.20

m1 n3 a1 vss vss n w=34u l=2u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
m2 z b vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m3 n1 a2 vdd vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
m4 z c n2 vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
m5 z a2 n3 vss n w=34u l=2u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
m6 n1 a1 vdd vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
m7 z c vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m8 n2 b n1 vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
.ends
