* Mon Aug 16 14:10:59 CEST 2004
.subckt nd2v0x8 a b vdd vss z 
*SPICE circuit <nd2v0x8> from XCircuit v3.10

m1 n1 a vss vss n w=80u l=2.3636u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m2 z a vdd vdd p w=96u l=2.3636u ad='96u*5u+12p' as='96u*5u+12p' pd='96u*2+14u' ps='96u*2+14u'
m3 z b n1 vss n w=80u l=2.3636u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m4 z b vdd vdd p w=96u l=2.3636u ad='96u*5u+12p' as='96u*5u+12p' pd='96u*2+14u' ps='96u*2+14u'
.ends
