magic
tech scmos
timestamp 1522931348
<< pwell >>
rect 0 0 152 36
rect 2 -3 72 0
<< nwell >>
rect 0 36 152 80
<< polysilicon >>
rect 13 70 15 74
rect 59 72 115 74
rect 59 64 61 72
rect 69 64 71 68
rect 79 64 81 68
rect 86 64 88 72
rect 96 64 98 68
rect 103 64 105 68
rect 23 56 25 61
rect 42 58 44 63
rect 49 58 51 63
rect 13 38 15 42
rect 23 39 25 42
rect 23 38 38 39
rect 13 37 19 38
rect 23 37 33 38
rect 13 33 14 37
rect 18 33 19 37
rect 13 32 19 33
rect 31 34 33 37
rect 37 34 38 38
rect 31 33 38 34
rect 13 28 15 32
rect 31 30 33 33
rect 42 23 44 52
rect 49 48 51 52
rect 49 47 55 48
rect 49 43 50 47
rect 54 43 55 47
rect 49 42 55 43
rect 59 38 61 52
rect 49 36 61 38
rect 49 23 51 36
rect 69 33 71 52
rect 79 48 81 58
rect 75 47 81 48
rect 75 43 76 47
rect 80 43 81 47
rect 75 42 81 43
rect 69 32 75 33
rect 55 31 61 32
rect 55 27 56 31
rect 60 27 61 31
rect 55 26 61 27
rect 59 23 61 26
rect 69 28 70 32
rect 74 28 75 32
rect 69 27 75 28
rect 69 23 71 27
rect 79 23 81 42
rect 86 38 88 58
rect 113 62 115 72
rect 133 63 135 68
rect 96 48 98 51
rect 92 47 98 48
rect 92 43 93 47
rect 97 43 98 47
rect 92 42 98 43
rect 103 39 105 51
rect 113 48 115 51
rect 133 49 135 53
rect 126 48 135 49
rect 113 46 121 48
rect 119 39 121 46
rect 126 44 127 48
rect 131 44 135 48
rect 126 43 135 44
rect 103 38 109 39
rect 86 36 98 38
rect 86 31 92 32
rect 86 27 87 31
rect 91 27 92 31
rect 86 26 92 27
rect 86 23 88 26
rect 96 23 98 36
rect 103 34 104 38
rect 108 34 109 38
rect 103 33 109 34
rect 119 38 125 39
rect 119 34 120 38
rect 124 34 125 38
rect 119 33 125 34
rect 103 23 105 33
rect 123 30 125 33
rect 133 30 135 43
rect 31 18 33 23
rect 123 19 125 24
rect 133 18 135 23
rect 13 11 15 14
rect 42 11 44 17
rect 49 12 51 17
rect 13 9 44 11
rect 38 6 40 9
rect 59 8 61 17
rect 69 12 71 17
rect 79 12 81 17
rect 86 8 88 17
rect 96 12 98 17
rect 103 12 105 17
rect 59 6 88 8
rect 38 4 49 6
rect 47 -9 49 4
<< ndiffusion >>
rect 24 29 31 30
rect 6 27 13 28
rect 6 23 7 27
rect 11 23 13 27
rect 6 22 13 23
rect 8 14 13 22
rect 15 20 20 28
rect 24 25 25 29
rect 29 25 31 29
rect 24 24 31 25
rect 26 23 31 24
rect 33 23 40 30
rect 116 29 123 30
rect 116 25 117 29
rect 121 25 123 29
rect 116 24 123 25
rect 125 29 133 30
rect 125 25 127 29
rect 131 25 133 29
rect 125 24 133 25
rect 15 19 22 20
rect 15 15 17 19
rect 21 15 22 19
rect 35 22 42 23
rect 35 18 36 22
rect 40 18 42 22
rect 35 17 42 18
rect 44 17 49 23
rect 51 22 59 23
rect 51 18 53 22
rect 57 18 59 22
rect 51 17 59 18
rect 61 22 69 23
rect 61 18 63 22
rect 67 18 69 22
rect 61 17 69 18
rect 71 22 79 23
rect 71 18 73 22
rect 77 18 79 22
rect 71 17 79 18
rect 81 17 86 23
rect 88 22 96 23
rect 88 18 90 22
rect 94 18 96 22
rect 88 17 96 18
rect 98 17 103 23
rect 105 22 112 23
rect 105 18 107 22
rect 111 18 112 22
rect 127 23 133 24
rect 135 29 142 30
rect 135 25 137 29
rect 141 25 142 29
rect 135 23 142 25
rect 105 17 112 18
rect 15 14 22 15
<< pdiffusion >>
rect 8 56 13 70
rect 6 54 13 56
rect 6 50 7 54
rect 11 50 13 54
rect 6 47 13 50
rect 6 43 7 47
rect 11 43 13 47
rect 6 42 13 43
rect 15 69 22 70
rect 15 65 17 69
rect 21 65 22 69
rect 15 64 22 65
rect 15 56 21 64
rect 54 58 59 64
rect 34 57 42 58
rect 15 55 23 56
rect 15 51 17 55
rect 21 51 23 55
rect 15 42 23 51
rect 25 48 30 56
rect 34 53 35 57
rect 39 53 42 57
rect 34 52 42 53
rect 44 52 49 58
rect 51 57 59 58
rect 51 53 53 57
rect 57 53 59 57
rect 51 52 59 53
rect 61 57 69 64
rect 61 53 63 57
rect 67 53 69 57
rect 61 52 69 53
rect 71 63 79 64
rect 71 59 73 63
rect 77 59 79 63
rect 71 58 79 59
rect 81 58 86 64
rect 88 63 96 64
rect 88 59 90 63
rect 94 59 96 63
rect 88 58 96 59
rect 71 52 77 58
rect 25 47 32 48
rect 25 43 27 47
rect 31 43 32 47
rect 25 42 32 43
rect 91 51 96 58
rect 98 51 103 64
rect 105 62 110 64
rect 126 62 133 63
rect 105 61 113 62
rect 105 57 107 61
rect 111 57 113 61
rect 105 51 113 57
rect 115 57 120 62
rect 126 58 127 62
rect 131 58 133 62
rect 115 56 122 57
rect 115 52 117 56
rect 121 52 122 56
rect 126 53 133 58
rect 135 59 140 63
rect 135 58 142 59
rect 135 54 137 58
rect 141 54 142 58
rect 135 53 142 54
rect 115 51 122 52
<< metal1 >>
rect 2 72 150 76
rect 2 69 31 72
rect 2 68 17 69
rect 21 68 31 69
rect 35 68 41 72
rect 45 68 122 72
rect 126 68 150 72
rect 17 55 21 65
rect 6 54 11 55
rect 6 50 7 54
rect 35 57 39 68
rect 73 63 77 68
rect 73 58 77 59
rect 85 59 90 63
rect 94 59 95 63
rect 106 61 112 68
rect 63 57 67 58
rect 35 52 39 53
rect 42 53 53 57
rect 57 53 58 57
rect 17 50 21 51
rect 6 47 11 50
rect 6 43 7 47
rect 11 43 19 46
rect 6 42 19 43
rect 25 43 27 47
rect 31 43 32 47
rect 6 28 10 42
rect 25 37 29 43
rect 42 38 46 53
rect 63 47 67 53
rect 49 43 50 47
rect 13 33 14 37
rect 18 33 29 37
rect 32 34 33 38
rect 37 34 48 38
rect 25 29 29 33
rect 6 27 11 28
rect 6 23 7 27
rect 25 24 29 25
rect 6 22 11 23
rect 36 22 40 23
rect 17 19 21 20
rect 17 12 21 15
rect 44 22 48 34
rect 54 32 58 47
rect 63 43 76 47
rect 80 43 81 47
rect 54 31 60 32
rect 54 27 56 31
rect 54 26 60 27
rect 63 22 67 43
rect 85 40 89 59
rect 106 57 107 61
rect 111 57 112 61
rect 126 62 132 68
rect 126 58 127 62
rect 131 58 132 62
rect 137 58 141 59
rect 117 56 121 57
rect 80 36 89 40
rect 93 52 117 54
rect 93 50 121 52
rect 93 47 97 50
rect 125 48 131 54
rect 125 46 127 48
rect 80 33 84 36
rect 70 32 84 33
rect 93 32 97 43
rect 101 38 107 46
rect 117 44 127 46
rect 117 42 131 44
rect 137 38 141 54
rect 101 34 104 38
rect 108 34 111 38
rect 119 34 120 38
rect 124 34 141 38
rect 74 28 84 32
rect 70 27 84 28
rect 44 18 53 22
rect 57 18 58 22
rect 36 12 40 18
rect 63 17 67 18
rect 73 22 77 23
rect 80 22 84 27
rect 87 31 97 32
rect 91 30 97 31
rect 91 29 122 30
rect 91 27 117 29
rect 87 26 117 27
rect 116 25 117 26
rect 121 25 122 29
rect 127 29 131 30
rect 80 18 90 22
rect 94 18 95 22
rect 106 18 107 22
rect 111 18 112 22
rect 73 12 77 18
rect 106 12 112 18
rect 127 12 131 25
rect 137 29 141 34
rect 137 24 141 25
rect 2 8 123 12
rect 127 8 134 12
rect 138 8 150 12
rect 2 4 150 8
rect 2 -3 72 4
rect 16 -22 22 -14
<< metal2 >>
rect 111 -20 114 33
rect 66 -23 114 -20
<< ntransistor >>
rect 13 14 15 28
rect 31 23 33 30
rect 123 24 125 30
rect 42 17 44 23
rect 49 17 51 23
rect 59 17 61 23
rect 69 17 71 23
rect 79 17 81 23
rect 86 17 88 23
rect 96 17 98 23
rect 103 17 105 23
rect 133 23 135 30
<< ptransistor >>
rect 13 42 15 70
rect 23 42 25 56
rect 42 52 44 58
rect 49 52 51 58
rect 59 52 61 64
rect 69 52 71 64
rect 79 58 81 64
rect 86 58 88 64
rect 96 51 98 64
rect 103 51 105 64
rect 113 51 115 62
rect 133 53 135 63
<< polycontact >>
rect 14 33 18 37
rect 33 34 37 38
rect 50 43 54 47
rect 76 43 80 47
rect 56 27 60 31
rect 70 28 74 32
rect 93 43 97 47
rect 127 44 131 48
rect 87 27 91 31
rect 104 34 108 38
rect 120 34 124 38
<< ndcontact >>
rect 7 23 11 27
rect 25 25 29 29
rect 117 25 121 29
rect 127 25 131 29
rect 17 15 21 19
rect 36 18 40 22
rect 53 18 57 22
rect 63 18 67 22
rect 73 18 77 22
rect 90 18 94 22
rect 107 18 111 22
rect 137 25 141 29
<< pdcontact >>
rect 7 50 11 54
rect 7 43 11 47
rect 17 65 21 69
rect 17 51 21 55
rect 35 53 39 57
rect 53 53 57 57
rect 63 53 67 57
rect 73 59 77 63
rect 90 59 94 63
rect 27 43 31 47
rect 107 57 111 61
rect 127 58 131 62
rect 117 52 121 56
rect 137 54 141 58
<< m2contact >>
rect 111 33 115 37
rect 62 -23 66 -19
<< psubstratepcontact >>
rect 123 8 127 12
rect 134 8 138 12
<< nsubstratencontact >>
rect 31 68 35 72
rect 41 68 45 72
rect 122 68 126 72
<< psubstratepdiff >>
rect 116 12 145 13
rect 116 8 123 12
rect 127 8 134 12
rect 138 8 145 12
rect 116 7 145 8
<< nsubstratendiff >>
rect 26 72 50 73
rect 26 68 31 72
rect 35 68 41 72
rect 45 68 50 72
rect 26 67 50 68
rect 121 72 127 73
rect 121 68 122 72
rect 126 68 127 72
rect 121 67 127 68
use ../pharosc_8.4/magic/cells/vsclib/mxn2v0x05  mxn2v0x05_0
timestamp 1522931348
transform -1 0 68 0 -1 0
box -4 -4 68 76
<< labels >>
rlabel polycontact 16 35 16 35 6 zn
rlabel polycontact 34 36 34 36 6 n4
rlabel polycontact 58 29 58 29 6 ci
rlabel polycontact 52 45 52 45 6 ci
rlabel polycontact 72 30 72 30 6 n1
rlabel polycontact 89 29 89 29 6 ci
rlabel polycontact 95 45 95 45 6 ci
rlabel polycontact 78 45 78 45 6 n2
rlabel polycontact 122 36 122 36 6 cn
rlabel metal1 21 35 21 35 6 zn
rlabel metal1 8 40 8 40 6 z
rlabel metal1 16 44 16 44 6 z
rlabel metal1 27 35 27 35 6 zn
rlabel metal1 51 20 51 20 6 n4
rlabel polycontact 57 29 57 29 6 ci
rlabel metal1 40 36 40 36 6 n4
rlabel polycontact 53 45 53 45 6 ci
rlabel metal1 50 55 50 55 6 n4
rlabel metal1 76 8 76 8 6 vss
rlabel metal1 77 30 77 30 6 n1
rlabel metal1 72 45 72 45 6 n2
rlabel metal1 65 37 65 37 6 n2
rlabel metal1 76 72 76 72 6 vdd
rlabel metal1 87 20 87 20 6 n1
rlabel metal1 104 40 104 40 6 d
rlabel metal1 95 40 95 40 6 ci
rlabel metal1 90 61 90 61 6 n1
rlabel metal1 104 28 104 28 6 ci
rlabel metal1 130 36 130 36 6 cn
rlabel metal1 120 44 120 44 6 cp
rlabel metal1 128 48 128 48 6 cp
rlabel metal1 139 41 139 41 6 cn
rlabel pdcontact 119 53 119 53 6 ci
<< end >>
