magic
tech scmos
timestamp 1523081934
<< metal1 >>
rect 271 231 311 236
rect 573 235 652 238
rect 627 221 631 229
rect 262 157 299 162
rect 262 156 302 157
rect 624 81 626 85
rect 271 74 311 80
rect 620 76 626 78
rect 624 74 626 76
rect 271 11 301 12
rect 271 7 299 11
rect 271 4 301 7
rect 553 5 652 10
<< metal2 >>
rect 692 232 716 236
rect 284 195 290 199
rect 349 200 358 204
rect 354 199 358 200
rect 393 199 397 205
rect 671 158 684 161
rect 330 127 334 131
rect 279 119 287 124
rect 619 95 628 99
rect 624 93 628 95
rect 608 81 620 85
rect 705 77 716 81
rect 602 75 620 76
rect 608 72 620 75
rect 317 54 320 55
rect 319 48 320 54
rect 317 47 320 48
rect 279 41 283 47
rect 659 7 665 11
rect 613 -52 627 -48
<< metal3 >>
rect 289 205 328 206
rect 289 201 322 205
rect 289 194 290 201
rect 297 200 322 201
rect 327 200 328 205
rect 297 199 328 200
rect 343 205 350 251
rect 715 236 723 237
rect 715 230 716 236
rect 722 230 723 236
rect 343 200 344 205
rect 349 200 350 205
rect 343 199 350 200
rect 369 215 619 222
rect 297 194 298 199
rect 289 193 298 194
rect 322 194 328 199
rect 369 194 376 215
rect 322 188 376 194
rect 286 125 296 126
rect 286 119 287 125
rect 293 120 532 125
rect 293 119 608 120
rect 286 118 296 119
rect 526 114 608 119
rect 602 88 608 114
rect 612 101 619 215
rect 664 161 672 162
rect 664 155 665 161
rect 671 155 672 161
rect 612 100 620 101
rect 612 94 613 100
rect 619 94 620 100
rect 612 93 620 94
rect 601 87 609 88
rect 601 81 602 87
rect 608 81 609 87
rect 601 80 609 81
rect 601 75 609 76
rect 601 69 602 75
rect 608 69 609 75
rect 278 54 320 55
rect 278 52 313 54
rect 278 47 279 52
rect 284 48 313 52
rect 319 48 320 54
rect 601 50 609 69
rect 284 47 320 48
rect 278 46 320 47
rect 342 46 609 50
rect 342 41 343 46
rect 348 44 609 46
rect 348 41 349 44
rect 601 43 609 44
rect 342 40 349 41
rect 664 12 672 155
rect 715 82 723 230
rect 715 76 716 82
rect 722 76 723 82
rect 715 75 723 76
rect 664 6 665 12
rect 671 6 672 12
rect 664 5 672 6
<< m2contact >>
rect 688 232 692 236
rect 354 195 358 199
rect 393 195 397 199
rect 299 157 303 162
rect 684 158 688 162
rect 330 123 334 127
rect 624 89 628 93
rect 620 81 624 85
rect 701 77 705 81
rect 620 72 624 76
rect 299 7 303 11
rect 655 7 659 11
rect 609 -52 613 -48
<< m3contact >>
rect 716 230 722 236
rect 290 194 297 201
rect 322 200 327 205
rect 344 200 349 205
rect 665 155 671 161
rect 287 119 293 125
rect 613 94 619 100
rect 602 81 608 87
rect 716 76 722 82
rect 602 69 608 75
rect 279 47 284 52
rect 313 48 319 54
rect 343 41 348 46
rect 665 6 671 12
use ./decoder  decoder_0
timestamp 1523081934
transform 1 0 58 0 1 160
box -58 -160 229 80
use ./comp  comp_0
timestamp 1523081934
transform 1 0 323 0 1 160
box -22 -240 296 83
use 3_bitmux  3_bitmux_0
timestamp 1523081934
transform 1 0 654 0 1 160
box -29 -160 85 80
<< labels >>
rlabel metal2 331 129 331 129 1 e
rlabel metal2 396 200 396 200 1 f
rlabel metal3 346 246 346 246 5 d
rlabel metal2 625 -50 625 -50 7 out
rlabel metal1 629 228 629 228 1 sel
<< end >>
