* Spice description of vfeed2
* Spice driver version 134999461
* Date 31/05/2007 at 21:35:58
* vxlib 0.13um values
.subckt vfeed2 vdd vss
.ends
