* Thu Jan 27 22:08:43 CET 2005
.subckt nr2v0x6 a b vdd vss z 
*SPICE circuit <nr2v0x6> from XCircuit v3.10

m1 z a vss vss n w=45u l=2u ad='45u*5u+12p' as='45u*5u+12p' pd='45u*2+14u' ps='45u*2+14u'
m2 n1 a vdd vdd p w=168u l=2u ad='168u*5u+12p' as='168u*5u+12p' pd='168u*2+14u' ps='168u*2+14u'
m3 z b vss vss n w=45u l=2u ad='45u*5u+12p' as='45u*5u+12p' pd='45u*2+14u' ps='45u*2+14u'
m4 z b n1 vdd p w=168u l=2u ad='168u*5u+12p' as='168u*5u+12p' pd='168u*2+14u' ps='168u*2+14u'
.ends
