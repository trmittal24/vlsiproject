* Spice description of iv1_x3
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:09
*
.subckt iv1_x3 a vdd vss z 
M2  vdd   a     z     vdd p  L=0.13U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U  
M1  z     a     vdd   vdd p  L=0.13U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U  
M4  z     a     vss   vss n  L=0.13U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U  
M3  vss   a     z     vss n  L=0.13U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U  
C4  a     vss   1.313f
C3  vdd   vss   1.468f
C2  z     vss   2.307f
.ends
