* Spice description of iv1_x05
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:09
*
.subckt iv1_x05 a vdd vss z 
M1  vdd   a     z     vdd p  L=0.13U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U  
M2  vss   a     z     vss n  L=0.13U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U  
C4  a     vss   0.736f
C3  vdd   vss   0.917f
C1  z     vss   1.391f
.ends
