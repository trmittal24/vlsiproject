* Wed Apr 11 10:41:37 CEST 2007
.subckt xor2v0x3 a b vdd vss z
*SPICE circuit <xor2v0x3> from XCircuit v3.4 rev 26

m1 z bn an vdd p w=54u l=2u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m2 bn b vss vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m3 an a vss vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m4 z an n1 vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m5 n1 bn vss vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m6 an a vdd vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m7 bn b vdd vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m8 z b an vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m9 z an bn vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
.ends
