* Tue Aug 10 11:21:06 CEST 2004
.subckt aoi21_x2 a1 a2 b vdd vss z 
*SPICE circuit <aoi21_x2> from XCircuit v3.10

m1 n1 a2 vdd vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
m2 n1 a1 vdd vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
m3 n2 a1 vss vss n w=33u l=2.3636u ad='33u*5u+12p' as='33u*5u+12p' pd='33u*2+14u' ps='33u*2+14u'
m4 z b vss vss n w=22u l=2.3636u ad='22u*5u+12p' as='22u*5u+12p' pd='22u*2+14u' ps='22u*2+14u'
m5 z a2 n2 vss n w=33u l=2.3636u ad='33u*5u+12p' as='33u*5u+12p' pd='33u*2+14u' ps='33u*2+14u'
m6 z b n1 vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
.ends
