magic
tech scmos
timestamp 1522414328
<< metal1 >>
rect 706 -318 785 -314
rect 706 -400 710 -318
rect 1005 -327 1266 -323
rect 724 -341 792 -338
rect 724 -390 727 -341
rect 827 -363 831 -349
rect 785 -366 831 -363
rect 836 -389 840 -347
rect 940 -349 951 -348
rect 940 -352 948 -349
rect 762 -390 840 -389
rect 766 -392 840 -390
rect 932 -390 935 -352
rect 1012 -391 1015 -377
rect 1030 -388 1049 -385
rect 723 -401 769 -398
rect 984 -401 1030 -398
rect 1263 -482 1266 -327
rect 665 -587 668 -564
rect 688 -588 701 -585
rect 627 -613 631 -608
rect 698 -623 701 -588
rect 888 -612 892 -608
rect 674 -627 701 -623
rect 940 -656 1019 -653
rect 752 -663 763 -660
<< metal2 >>
rect 781 -383 784 -366
rect 690 -385 784 -383
rect 507 -386 784 -385
rect 793 -383 796 -350
rect 845 -374 849 -346
rect 952 -353 1040 -350
rect 845 -377 1012 -374
rect 793 -384 1030 -383
rect 793 -386 1026 -384
rect 507 -388 693 -386
rect 507 -598 510 -388
rect 762 -448 765 -394
rect 1012 -445 1015 -395
rect 1037 -396 1040 -353
rect 1053 -388 1272 -385
rect 1012 -448 1044 -445
rect 762 -451 784 -448
rect 763 -481 773 -478
rect 781 -495 784 -451
rect 1023 -482 1033 -479
rect 1041 -492 1044 -448
rect 767 -498 784 -495
rect 1027 -495 1044 -492
rect 753 -514 759 -511
rect 622 -660 625 -613
rect 622 -663 748 -660
rect 756 -669 759 -514
rect 767 -598 770 -498
rect 948 -588 957 -583
rect 884 -653 887 -612
rect 884 -656 936 -653
rect 944 -660 947 -606
rect 767 -663 947 -660
rect 954 -669 957 -588
rect 756 -672 957 -669
rect 1010 -669 1013 -514
rect 1027 -598 1030 -495
rect 1269 -510 1272 -388
rect 1209 -588 1216 -584
rect 1020 -660 1023 -656
rect 1203 -660 1206 -607
rect 1020 -663 1206 -660
rect 1213 -669 1216 -588
rect 1010 -672 1216 -669
<< m2contact >>
rect 781 -366 785 -362
rect 724 -394 728 -390
rect 762 -394 766 -390
rect 948 -353 952 -349
rect 1012 -377 1016 -373
rect 932 -394 936 -390
rect 1026 -388 1030 -384
rect 1049 -388 1053 -384
rect 1012 -395 1016 -391
rect 759 -482 763 -478
rect 773 -482 777 -478
rect 1019 -482 1023 -478
rect 1033 -482 1037 -478
rect 749 -514 753 -510
rect 1009 -514 1013 -510
rect 1269 -514 1273 -510
rect 622 -613 627 -608
rect 884 -612 888 -608
rect 936 -656 940 -652
rect 1019 -656 1023 -652
rect 748 -663 752 -659
rect 763 -663 767 -659
use mux  mux_0
timestamp 1522414328
transform 0 -1 857 1 0 -323
box -29 -160 85 80
use diff2  diff2_0
timestamp 1522414328
transform 1 0 511 0 1 -473
box -4 -160 252 80
use diff2  diff2_1
timestamp 1522414328
transform 1 0 771 0 1 -473
box -4 -160 252 80
use diff2  diff2_2
timestamp 1522414328
transform 1 0 1031 0 1 -473
box -4 -160 252 80
<< end >>
