* Tue Aug 10 11:21:07 CEST 2004
.subckt iv1_x4 a vdd vss z 
*SPICE circuit <iv1_x4> from XCircuit v3.10

m1 z a vss vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m2 z a vdd vdd p w=76u l=2u ad='76u*5u+12p' as='76u*5u+12p' pd='76u*2+14u' ps='76u*2+14u'
.ends
