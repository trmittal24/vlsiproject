* Spice description of oai21a2bv0x05
* Spice driver version 134999461
* Date 17/05/2007 at  9:29:37
* wsclib 0.13um values
.subckt oai21a2bv0x05 a1 a2 b vdd vss z
M01 vdd   a1    01    vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M02 04    a1    vss   vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M03 01    a2n   z     vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M04 vss   a2n   04    vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M05 z     bn    vdd   vdd p  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M06 04    bn    z     vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M07 bn    b     vdd   vdd p  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
M08 vdd   a2    a2n   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M09 bn    b     vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M10 vss   a2    a2n   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
C6  04    vss   0.231f
C8  a1    vss   0.397f
C5  a2    vss   0.368f
C3  a2n   vss   0.954f
C4  b     vss   0.399f
C1  bn    vss   0.517f
C7  z     vss   0.591f
.ends
