* Mon Aug 16 14:22:56 CEST 2004
.subckt inv_x8 i nq vdd vss 
*SPICE circuit <inv_x8> from XCircuit v3.10

m1 nq i vss vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m2 nq i vdd vdd p w=160u l=2u ad='160u*5u+12p' as='160u*5u+12p' pd='160u*2+14u' ps='160u*2+14u'
.ends
