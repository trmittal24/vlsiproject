* Sun Apr  2 13:48:00 CEST 2006
.subckt or2v0x05 a b vdd vss z 
*SPICE circuit <or2v0x05> from XCircuit v3.20

m1 z zn vdd vdd p w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m2 z zn vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m3 zn a vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m4 n1 a vdd vdd p w=17u l=2u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m5 zn b vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m6 zn b n1 vdd p w=17u l=2u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
.ends
