* Spice description of na4_x4
* Spice driver version 134999461
* Date 31/05/2007 at 10:38:08
* ssxlib 0.13um values
.subckt na4_x4 i0 i1 i2 i3 nq vdd vss
Mtr_00001 sig3  sig4  vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00002 vss   sig3  nq    vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00003 nq    sig3  vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00004 sig8  i3    sig4  vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00005 vss   i0    sig5  vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00006 sig5  i1    sig9  vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00007 sig9  i2    sig8  vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00008 vdd   sig4  sig3  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00009 vdd   sig3  nq    vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
Mtr_00010 nq    sig3  vdd   vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
Mtr_00011 sig4  i0    vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00012 vdd   i1    sig4  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00013 sig4  i2    vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00014 vdd   i3    sig4  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
C6  i0    vss   0.768f
C7  i1    vss   0.790f
C11 i2    vss   0.813f
C10 i3    vss   0.827f
C2  nq    vss   0.645f
C3  sig3  vss   0.794f
C4  sig4  vss   1.367f
.ends
