* Spice description of vddtie
* Spice driver version 134999461
* Date  6/02/2007 at 12:03:55
* rgalib 0.13um values
.subckt vddtie vdd vss z
Mtr_00001 z     vss   sig2  vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00002 sig3  vss   z     vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00003 z     vss   vdd   vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
Mtr_00004 vdd   vss   z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
C1  z     vss   0.660f
.ends
