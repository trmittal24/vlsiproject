* Sun Apr  2 13:48:07 CEST 2006
.subckt or2v0x4 a b vdd vss z 
*SPICE circuit <or2v0x4> from XCircuit v3.20

m1 z zn vdd vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m2 z zn vss vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m3 zn a vss vss n w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m4 n1 a vdd vdd p w=42u l=2u ad='42u*5u+12p' as='42u*5u+12p' pd='42u*2+14u' ps='42u*2+14u'
m5 zn b vss vss n w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m6 zn b n1 vdd p w=42u l=2u ad='42u*5u+12p' as='42u*5u+12p' pd='42u*2+14u' ps='42u*2+14u'
.ends
