* Spice description of nao2o22_x1
* Spice driver version 134999461
* Date 31/05/2007 at 10:38:14
* ssxlib 0.13um values
.subckt nao2o22_x1 i0 i1 i2 i3 nq vdd vss
Mtr_00001 vss   i2    sig2  vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00002 sig2  i3    vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00003 nq    i1    sig2  vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00004 sig2  i0    nq    vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00005 nq    i1    sig8  vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
Mtr_00006 sig8  i0    vdd   vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
Mtr_00007 sig10 i3    nq    vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
Mtr_00008 vdd   i2    sig10 vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
C4  i0    vss   0.624f
C3  i1    vss   0.652f
C6  i2    vss   0.732f
C7  i3    vss   0.759f
C1  nq    vss   0.776f
C2  sig2  vss   0.345f
.ends
