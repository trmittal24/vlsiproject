* Wed Apr  5 08:55:23 CEST 2006
.subckt bf1v2x8 a vdd vss z 
*SPICE circuit <bf1v2x8> from XCircuit v3.20

m1 an a vss vss n w=22u l=2.3636u ad='22u*5u+12p' as='22u*5u+12p' pd='22u*2+14u' ps='22u*2+14u'
m2 an a vdd vdd p w=44u l=2.3636u ad='44u*5u+12p' as='44u*5u+12p' pd='44u*2+14u' ps='44u*2+14u'
m3 z an vss vss n w=52u l=2.3636u ad='52u*5u+12p' as='52u*5u+12p' pd='52u*2+14u' ps='52u*2+14u'
m4 z an vdd vdd p w=104u l=2.3636u ad='104u*5u+12p' as='104u*5u+12p' pd='104u*2+14u' ps='104u*2+14u'
.ends
