magic
tech scmos
timestamp 1521311720
<< metal1 >>
rect 221 138 280 141
rect 474 133 523 136
rect 219 -8 223 74
rect 434 -7 438 71
rect 711 -7 717 68
rect 434 -8 719 -7
rect 219 -11 719 -8
<< metal2 >>
rect 336 30 340 42
rect 161 26 177 30
rect 336 27 370 30
rect 172 7 177 26
rect 367 7 370 27
rect 416 21 436 24
rect 172 3 370 7
rect 432 4 436 21
rect 601 23 604 40
rect 601 20 637 23
rect 633 4 637 20
rect 432 0 637 4
<< m2contact >>
rect 157 26 161 30
rect 412 21 416 25
use diff2  diff2_0
timestamp 1521310090
transform 1 0 8 0 1 70
box -8 -70 218 80
use diff2  diff2_1
timestamp 1521310090
transform 1 0 263 0 1 65
box -8 -70 218 80
use diff2  diff2_2
timestamp 1521310090
transform 1 0 527 0 1 62
box -8 -70 218 80
<< end >>
