* Spice description of inv_x2
* Spice driver version 134999461
* Date 21/07/2007 at 19:29:27
* sxlib 0.13um values
.subckt inv_x2 i nq vdd vss
Mtr_00001 vss   i     nq    vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00002 nq    i     vdd   vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
C4  i     vss   0.868f
C1  nq    vss   0.906f
.ends
