* Wed Apr  5 08:58:30 CEST 2006
.subckt bf1v0x8 a vdd vss z 
*SPICE circuit <bf1v0x8> from XCircuit v3.20

m1 an a vss vss n w=23u l=2u ad='23u*5u+12p' as='23u*5u+12p' pd='23u*2+14u' ps='23u*2+14u'
m2 an a vdd vdd p w=43u l=2u ad='43u*5u+12p' as='43u*5u+12p' pd='43u*2+14u' ps='43u*2+14u'
m3 z an vss vss n w=52u l=2u ad='52u*5u+12p' as='52u*5u+12p' pd='52u*2+14u' ps='52u*2+14u'
m4 z an vdd vdd p w=104u l=2u ad='104u*5u+12p' as='104u*5u+12p' pd='104u*2+14u' ps='104u*2+14u'
.ends
