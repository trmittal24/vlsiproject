* Spice description of an2_x05
* Spice driver version 134999461
* Date 31/05/2007 at 21:32:09
* vxlib 0.13um values
.subckt an2_x05 a b vdd vss z
M1a vdd   a     zn    vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M1b zn    b     vdd   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M1z z     zn    vdd   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M2a n1    a     vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
M2b zn    b     n1    vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
M2z vss   zn    z     vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
C6  a     vss   0.561f
C7  b     vss   0.638f
C3  z     vss   0.663f
C4  zn    vss   0.704f
.ends
