* Spice description of iv1v7x1
* Spice driver version 134999461
* Date 17/05/2007 at  9:14:04
* vsclib 0.13um values
.subckt iv1v7x1 a vdd vss z
M01 z     a     vdd   vdd p  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
M02 vss   a     z     vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
C3  a     vss   0.498f
C2  z     vss   0.412f
.ends
