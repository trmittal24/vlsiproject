* Mon Aug 16 14:10:57 CEST 2004
.subckt aoi22v0x2 a1 a2 b1 b2 vdd vss z 
*SPICE circuit <aoi22v0x2> from XCircuit v3.10

m1 n1 b1 vss vss n w=25u l=2.3636u ad='25u*5u+12p' as='25u*5u+12p' pd='25u*2+14u' ps='25u*2+14u'
m2 z b1 n3 vdd p w=56u l=2.3636u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m3 n3 a1 vdd vdd p w=56u l=2.3636u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m4 n3 a2 vdd vdd p w=56u l=2.3636u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m5 n2 a1 vss vss n w=25u l=2.3636u ad='25u*5u+12p' as='25u*5u+12p' pd='25u*2+14u' ps='25u*2+14u'
m6 z b2 n1 vss n w=25u l=2.3636u ad='25u*5u+12p' as='25u*5u+12p' pd='25u*2+14u' ps='25u*2+14u'
m7 z a2 n2 vss n w=25u l=2.3636u ad='25u*5u+12p' as='25u*5u+12p' pd='25u*2+14u' ps='25u*2+14u'
m8 z b2 n3 vdd p w=56u l=2.3636u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
.ends
