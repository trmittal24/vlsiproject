* Thu Jan 11 12:50:31 CET 2007
.subckt mxi2v0x1 a0 a1 s vdd vss z
