* Sat Aug 27 19:34:36 CEST 2005
.subckt nd2v4x8 a b vdd vss z 
*SPICE circuit <nd2v4x8> from XCircuit v3.20

m1 n1 a vss vss n w=52u l=2.3636u ad='52u*5u+12p' as='52u*5u+12p' pd='52u*2+14u' ps='52u*2+14u'
m2 z a vdd vdd p w=125u l=2.3636u ad='125u*5u+12p' as='125u*5u+12p' pd='125u*2+14u' ps='125u*2+14u'
m3 z b n1 vss n w=52u l=2.3636u ad='52u*5u+12p' as='52u*5u+12p' pd='52u*2+14u' ps='52u*2+14u'
m4 z b vdd vdd p w=125u l=2.3636u ad='125u*5u+12p' as='125u*5u+12p' pd='125u*2+14u' ps='125u*2+14u'
.ends
