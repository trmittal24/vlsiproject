* Sat Aug 27 22:10:25 CEST 2005
.subckt iv1v5x2 a vdd vss z 
*SPICE circuit <iv1v5x2> from XCircuit v3.20

m1 z a vss vss n w=11u l=2u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m2 z a vdd vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
.ends
