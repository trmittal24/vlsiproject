* Thu Sep  1 18:58:50 CEST 2005
.subckt nr2v1x6 a b vdd vss z 
*SPICE circuit <nr2v1x6> from XCircuit v3.20

m1 z a vss vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m2 n1 a vdd vdd p w=168u l=2u ad='168u*5u+12p' as='168u*5u+12p' pd='168u*2+14u' ps='168u*2+14u'
m3 z b vss vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m4 z b n1 vdd p w=168u l=2u ad='168u*5u+12p' as='168u*5u+12p' pd='168u*2+14u' ps='168u*2+14u'
.ends
