* Tue Aug 10 11:21:07 CEST 2004
.subckt oai22_x05 a1 a2 b1 b2 vdd vss z 
*SPICE circuit <oai22_x05> from XCircuit v3.10

m1 z b1 n2 vss n w=9u l=2u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m2 int14 b1 vdd vdd p w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m3 n1 a1 vdd vdd p w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m4 z b2 int14 vdd p w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m5 n2 a2 vss vss n w=9u l=2u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m6 n2 a1 vss vss n w=9u l=2u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m7 z b2 n2 vss n w=9u l=2u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m8 z a2 n1 vdd p w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
.ends
