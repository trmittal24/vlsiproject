magic
tech scmos
timestamp 1523173521
<< polysilicon >>
rect 832 -13 834 -4
rect 884 -217 886 -205
rect 901 -217 903 -205
rect 908 -217 910 -197
<< metal1 >>
rect 859 189 907 193
rect 857 104 898 108
rect 141 44 182 49
rect 177 -72 182 44
rect 858 26 883 29
rect 826 -18 829 -14
rect 177 -77 533 -72
rect 178 -78 533 -77
rect 31 -140 193 -134
rect 222 -140 277 -132
rect 218 -150 237 -147
rect 544 -161 548 -145
rect 544 -165 551 -161
rect 253 -201 256 -166
rect 572 -174 576 -149
rect 660 -159 820 -154
rect -11 -213 34 -202
rect 179 -212 227 -203
rect 884 -201 888 -196
rect 899 -201 903 -196
rect 908 -193 912 -188
rect 765 -220 851 -212
rect 729 -253 733 -246
rect 820 -262 844 -258
rect 766 -284 852 -276
rect 661 -325 666 -321
<< metal2 >>
rect 899 108 902 109
rect 395 44 439 49
rect 656 46 671 49
rect 435 -57 439 44
rect 73 -58 610 -57
rect 668 -58 671 46
rect 71 -60 673 -58
rect 71 -63 669 -60
rect 71 -166 75 -63
rect 267 -85 270 -84
rect 435 -85 439 -63
rect 604 -64 669 -63
rect 267 -88 439 -85
rect 267 -105 270 -88
rect 237 -108 270 -105
rect 237 -146 240 -108
rect 535 -146 539 -78
rect 241 -150 270 -147
rect 535 -149 572 -146
rect 267 -154 270 -150
rect 822 -153 826 -18
rect 205 -162 208 -157
rect 604 -158 655 -154
rect 205 -165 253 -162
rect 540 -163 565 -162
rect 535 -166 565 -163
rect 32 -169 75 -166
rect -39 -176 5 -173
rect -39 -251 -35 -176
rect 252 -238 255 -205
rect 734 -244 781 -242
rect 660 -245 777 -244
rect 660 -247 740 -245
rect -59 -255 -39 -251
rect 822 -321 826 -159
rect 884 -192 887 26
rect 899 -192 902 104
rect 908 -184 911 189
rect 884 -205 887 -196
rect 899 -205 902 -196
rect 908 -197 911 -188
rect 661 -325 828 -321
<< polycontact >>
rect 829 -18 834 -13
rect 908 -197 912 -193
rect 884 -205 888 -201
rect 899 -205 903 -201
<< m2contact >>
rect 907 189 911 193
rect 898 104 902 108
rect 883 26 887 30
rect 821 -18 826 -13
rect 669 -64 673 -60
rect 533 -78 539 -71
rect 237 -150 241 -146
rect 205 -157 209 -153
rect 267 -158 271 -154
rect 572 -149 577 -144
rect 28 -169 32 -165
rect 253 -166 257 -162
rect 5 -176 9 -172
rect 599 -159 604 -154
rect 655 -159 660 -154
rect 820 -159 826 -153
rect 908 -188 912 -184
rect 252 -205 256 -201
rect 884 -196 888 -192
rect 899 -196 903 -192
rect -39 -255 -35 -251
rect 777 -248 781 -244
rect 657 -325 661 -321
use totdiff3  totdiff3_0
timestamp 1523173042
transform 1 0 -552 0 1 620
box 507 -672 1412 -374
use bf1v0x4  bf1v0x4_0
timestamp 1523173042
transform -1 0 32 0 -1 -132
box -4 -4 44 76
use bf1v0x3  bf1v0x3_0
timestamp 1523173042
transform -1 0 223 0 -1 -132
box -4 -4 44 76
use 1counter  1counter_0
timestamp 1523173042
transform 1 0 544 0 1 -289
box -589 -79 227 161
use an2v0x3  an2v0x3_0
timestamp 1523173042
transform 1 0 775 0 1 -284
box -4 -4 60 76
use or3v0x3  or3v0x3_0
timestamp 1523173042
transform 1 0 839 0 1 -284
box -4 -4 84 76
<< labels >>
rlabel metal2 -57 -254 -57 -254 3 xxx
<< end >>
