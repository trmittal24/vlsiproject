* Mon Aug 16 14:10:57 CEST 2004
.subckt aoi21v0x2 a1 a2 b vdd vss z 
*SPICE circuit <aoi21v0x2> from XCircuit v3.10

m1 n1 a2 vdd vdd p w=54u l=2u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m2 n1 a1 vdd vdd p w=54u l=2u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m3 n2 a1 vss vss n w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m4 z b vss vss n w=15u l=2u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m5 z a2 n2 vss n w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m6 z b n1 vdd p w=54u l=2u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
.ends
