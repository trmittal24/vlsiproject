* Spice description of oa2a22_x2
* Spice driver version 134999461
* Date 31/05/2007 at 10:39:48
* ssxlib 0.13um values
.subckt oa2a22_x2 i0 i1 i2 i3 q vdd vss
Mtr_00001 sig3  i1    sig1  vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00002 vss   i0    sig3  vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00003 sig6  i3    vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00004 sig1  i2    sig6  vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00005 vss   sig1  q     vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00006 sig11 i1    sig1  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00007 sig11 i3    vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00008 vdd   i2    sig11 vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00009 sig1  i0    sig11 vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00010 q     sig1  vdd   vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
C4  i0    vss   0.660f
C5  i1    vss   0.688f
C7  i2    vss   0.688f
C8  i3    vss   0.660f
C9  q     vss   0.771f
C1  sig1  vss   0.994f
C11 sig11 vss   0.345f
.ends
