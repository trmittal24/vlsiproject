* Sat Aug 27 22:10:05 CEST 2005
.subckt iv1v4x4 a vdd vss z 
*SPICE circuit <iv1v4x4> from XCircuit v3.20

m1 z a vss vss n w=17u l=2u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m2 z a vdd vdd p w=68u l=2u ad='68u*5u+12p' as='68u*5u+12p' pd='68u*2+14u' ps='68u*2+14u'
.ends
