magic
tech scmos
timestamp 1523172170
<< metal1 >>
rect -34 228 56 236
rect 270 228 348 233
rect 286 195 330 199
rect 279 84 283 120
rect 317 88 324 92
rect 279 80 322 84
rect 304 53 308 80
rect 317 42 321 77
rect 285 38 321 42
rect 294 -199 299 38
rect 304 -192 308 21
rect 329 -49 333 92
rect 304 -196 319 -192
rect 294 -203 321 -199
rect -35 -274 59 -265
rect 272 -273 343 -268
<< metal2 >>
rect 72 231 76 235
rect 362 229 405 233
rect 287 185 324 189
rect 147 77 157 81
rect 208 6 238 10
rect 70 -47 76 -42
rect 287 -69 291 185
rect 287 -78 291 -74
rect 284 -82 291 -78
rect 295 176 323 180
rect 295 -96 299 176
rect 397 156 409 159
rect 362 79 380 83
rect 362 78 376 79
rect 304 25 308 49
rect 335 14 339 29
rect 311 10 339 14
rect 208 -118 220 -113
rect 295 -153 299 -101
rect 282 -157 299 -153
rect 311 -105 315 10
rect 384 5 409 8
rect 353 -47 357 -43
rect 320 -87 324 -74
rect 311 -109 323 -105
rect 154 -199 160 -193
rect 311 -235 315 -109
rect 404 -122 409 -118
rect 362 -197 376 -193
rect 362 -198 377 -197
rect 373 -201 377 -198
rect 282 -239 315 -235
rect 208 -271 239 -268
rect 383 -271 409 -268
rect 383 -272 412 -271
<< metal3 >>
rect 75 236 83 237
rect 75 230 76 236
rect 82 230 83 236
rect 75 88 83 230
rect 356 233 363 234
rect 356 229 357 233
rect 362 229 363 233
rect 201 162 209 163
rect 201 156 202 162
rect 208 156 209 162
rect 75 86 147 88
rect 75 84 148 86
rect 75 82 140 84
rect 75 -41 83 82
rect 139 77 140 82
rect 147 77 148 84
rect 139 76 148 77
rect 75 -47 76 -41
rect 82 -47 83 -41
rect 75 -191 83 -47
rect 201 11 209 156
rect 201 6 202 11
rect 208 6 209 11
rect 201 -112 209 6
rect 356 83 363 229
rect 356 78 357 83
rect 362 78 363 83
rect 356 -42 363 78
rect 356 -47 357 -42
rect 362 -47 363 -42
rect 285 -69 326 -68
rect 285 -74 286 -69
rect 291 -74 320 -69
rect 325 -74 326 -69
rect 285 -75 326 -74
rect 335 -95 342 -94
rect 294 -96 336 -95
rect 294 -101 295 -96
rect 300 -100 336 -96
rect 341 -100 342 -95
rect 300 -101 342 -100
rect 294 -102 335 -101
rect 201 -118 202 -112
rect 208 -118 209 -112
rect 75 -193 155 -191
rect 75 -197 147 -193
rect 146 -200 147 -197
rect 154 -200 155 -193
rect 146 -201 155 -200
rect 201 -266 209 -118
rect 356 -193 363 -47
rect 356 -198 357 -193
rect 362 -198 363 -193
rect 356 -199 363 -198
rect 408 159 415 160
rect 408 155 409 159
rect 414 155 415 159
rect 408 9 415 155
rect 408 5 409 9
rect 414 5 415 9
rect 408 -118 415 5
rect 408 -122 409 -118
rect 414 -122 415 -118
rect 201 -272 202 -266
rect 208 -272 209 -266
rect 408 -266 415 -122
rect 408 -271 409 -266
rect 414 -271 415 -266
rect 408 -272 415 -271
rect 201 -273 209 -272
<< m2contact >>
rect 67 231 72 236
rect 405 229 409 233
rect 393 156 397 160
rect 157 77 162 82
rect 304 49 308 53
rect 238 6 242 10
rect 65 -47 70 -42
rect 220 -118 225 -113
rect 160 -199 167 -192
rect 304 21 308 25
rect 376 75 380 79
rect 380 5 384 9
rect 349 -47 353 -43
rect 400 -122 404 -118
rect 377 -201 381 -197
rect 239 -271 243 -267
rect 379 -272 383 -268
<< m3contact >>
rect 76 230 82 236
rect 357 229 362 233
rect 202 156 208 162
rect 140 77 147 84
rect 202 6 208 11
rect 76 -47 82 -41
rect 286 -74 291 -69
rect 409 155 414 159
rect 357 78 362 83
rect 295 -101 300 -96
rect 202 -118 208 -112
rect 409 5 414 9
rect 357 -47 362 -42
rect 320 -74 325 -69
rect 336 -100 341 -95
rect 147 -200 154 -193
rect 409 -122 414 -118
rect 357 -198 362 -193
rect 202 -272 208 -266
rect 409 -271 414 -266
use decoder  decoder_0
timestamp 1523172170
transform 1 0 58 0 1 160
box -58 -160 229 80
use 3_bitmux  3_bitmux_0
timestamp 1523172170
transform 1 0 347 0 1 159
box -29 -160 85 80
use decoder  decoder_1
timestamp 1523172170
transform 1 0 58 0 1 -117
box -58 -160 229 80
use 3_bitmux  3_bitmux_1
timestamp 1523172170
transform 1 0 347 0 1 -117
box -29 -160 85 80
<< labels >>
rlabel metal1 -32 231 -32 231 3 vdd
rlabel metal1 -30 -270 -30 -270 3 gnd
<< end >>
