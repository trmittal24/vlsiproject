* Thu Sep  1 18:58:44 CEST 2005
.subckt nr2v1x2 a b vdd vss z 
*SPICE circuit <nr2v1x2> from XCircuit v3.20

m1 z a vss vss n w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m2 n1 a vdd vdd p w=54u l=2u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m3 z b vss vss n w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m4 z b n1 vdd p w=54u l=2u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
.ends
