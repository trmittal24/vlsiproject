* Tue Feb 20 08:57:11 CET 2007
.subckt nr2v0x2 a b vdd vss z
*SPICE circuit <nr2v0x2> from XCircuit v3.4 rev 26

m1 z a vss vss n w=36u l=2u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
m2 n1 a vdd vdd p w=52u l=2u ad='52u*5u+12p' as='52u*5u+12p' pd='52u*2+14u' ps='52u*2+14u'
m3 z b vss vss n w=36u l=2u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
m4 z b n1 vdd p w=52u l=2u ad='52u*5u+12p' as='52u*5u+12p' pd='52u*2+14u' ps='52u*2+14u'
.ends
