* Thu Jan 27 22:08:41 CET 2005
.subckt nr2v0x4 a b vdd vss z 
*SPICE circuit <nr2v0x4> from XCircuit v3.10

m1 z a vss vss n w=30u l=2.3636u ad='30u*5u+12p' as='30u*5u+12p' pd='30u*2+14u' ps='30u*2+14u'
m2 n1 a vdd vdd p w=112u l=2.3636u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
m3 z b vss vss n w=30u l=2.3636u ad='30u*5u+12p' as='30u*5u+12p' pd='30u*2+14u' ps='30u*2+14u'
m4 z b n1 vdd p w=112u l=2.3636u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
.ends
