* Mon Aug 16 14:22:56 CEST 2004
.subckt inv_x2 i nq vdd vss 
*SPICE circuit <inv_x2> from XCircuit v3.10

m1 nq i vss vss n w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m2 nq i vdd vdd p w=30u l=2.3636u ad='30u*5u+12p' as='30u*5u+12p' pd='30u*2+14u' ps='30u*2+14u'
.ends
