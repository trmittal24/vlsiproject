* Mon Aug 16 14:22:56 CEST 2004
.subckt inv_x1 i nq vdd vss 
*SPICE circuit <inv_x1> from XCircuit v3.10

m1 nq i vss vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m2 nq i vdd vdd p w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
.ends
