* Spice description of nd2_x2
* Spice driver version 134999461
* Date 31/05/2007 at 21:34:24
* vxlib 0.13um values
.subckt nd2_x2 a b vdd vss z
M1  z     b     vdd   vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M2  vdd   a     z     vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M3  z     b     n1    vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M4  n1    a     vss   vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
C6  a     vss   0.582f
C5  b     vss   0.450f
C3  z     vss   1.016f
.ends
