* Tue Dec 14 17:54:34 CET 2004
.subckt xnr3v1x1 a b c vdd vss z 
*SPICE circuit <xnr3v1x1> from XCircuit v3.20

m1 z cn izn vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m2 cn c vss vss n w=11u l=2u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m3 izn iz vss vss n w=13u l=2u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m4 n2 izn vss vss n w=13u l=2u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m5 z cn n2 vss n w=13u l=2u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m6 izn iz vdd vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m7 cn c vdd vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m8 z c izn vss n w=13u l=2u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m9 z izn cn vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m10 n1 bn vdd vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m11 iz b an vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m12 bn b vss vss n w=11u l=2u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m13 an a vss vss n w=11u l=2u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m14 iz an bn vss n w=14u l=2u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m15 an a vdd vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m16 bn b vdd vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m17 iz bn an vss n w=14u l=2u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m18 iz an n1 vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
.ends
