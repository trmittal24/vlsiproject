* Spice description of fulladder_x4
* Spice driver version 134999461
* Date 21/07/2007 at 19:29:14
* sxlib 0.13um values
.subckt fulladder_x4 a1 a2 a3 a4 b1 b2 b3 b4 cin1 cin2 cin3 cout sout vdd vss
Mtr_00001 vss   sig4  cout  vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00002 sig3  b2    vss   vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00003 vss   a2    sig3  vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00004 sig3  cin1  sig4  vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00005 sig1  a1    vss   vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00006 sig4  b1    sig1  vss n  L=0.12U  W=0.65U  AS=0.17225P  AD=0.17225P  PS=1.83U   PD=1.83U
Mtr_00007 cout  sig4  vss   vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00008 sout  sig15 vss   vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00009 vss   sig15 sout  vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00010 sig16 sig4  sig15 vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00011 vss   b4    sig16 vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00012 sig15 cin2  sig18 vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00013 sig18 b3    sig17 vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00014 sig16 a4    vss   vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00015 vss   cin3  sig16 vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00016 sig17 a3    vss   vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00017 cout  sig4  vdd   vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00018 sig6  b1    vdd   vdd p  L=0.12U  W=0.98U  AS=0.2597P   AD=0.2597P   PS=2.49U   PD=2.49U
Mtr_00019 sig4  cin1  sig6  vdd p  L=0.12U  W=0.98U  AS=0.2597P   AD=0.2597P   PS=2.49U   PD=2.49U
Mtr_00020 sig5  a2    sig4  vdd p  L=0.12U  W=1.42U  AS=0.3763P   AD=0.3763P   PS=3.37U   PD=3.37U
Mtr_00021 sig6  b2    sig5  vdd p  L=0.12U  W=1.42U  AS=0.3763P   AD=0.3763P   PS=3.37U   PD=3.37U
Mtr_00022 vdd   a1    sig6  vdd p  L=0.12U  W=0.98U  AS=0.2597P   AD=0.2597P   PS=2.49U   PD=2.49U
Mtr_00023 vdd   sig4  cout  vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00024 vdd   sig15 sout  vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00025 sout  sig15 vdd   vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00026 vdd   b3    sig25 vdd p  L=0.12U  W=0.76U  AS=0.2014P   AD=0.2014P   PS=2.05U   PD=2.05U
Mtr_00027 sig25 cin2  vdd   vdd p  L=0.12U  W=0.76U  AS=0.2014P   AD=0.2014P   PS=2.05U   PD=2.05U
Mtr_00028 sig25 b4    sig27 vdd p  L=0.12U  W=0.76U  AS=0.2014P   AD=0.2014P   PS=2.05U   PD=2.05U
Mtr_00029 sig27 a4    sig26 vdd p  L=0.12U  W=0.76U  AS=0.2014P   AD=0.2014P   PS=2.05U   PD=2.05U
Mtr_00030 sig25 a3    vdd   vdd p  L=0.12U  W=0.76U  AS=0.2014P   AD=0.2014P   PS=2.05U   PD=2.05U
Mtr_00031 sig15 sig4  sig25 vdd p  L=0.12U  W=0.98U  AS=0.2597P   AD=0.2597P   PS=2.49U   PD=2.49U
Mtr_00032 sig26 cin3  sig15 vdd p  L=0.12U  W=0.76U  AS=0.2014P   AD=0.2014P   PS=2.05U   PD=2.05U
C9  a1    vss   0.785f
C11 a2    vss   0.565f
C23 a3    vss   0.474f
C21 a4    vss   0.697f
C8  b1    vss   0.725f
C10 b2    vss   0.542f
C20 b3    vss   0.600f
C24 b4    vss   0.682f
C7  cin1  vss   0.652f
C19 cin2  vss   0.600f
C22 cin3  vss   0.586f
C13 cout  vss   0.734f
C15 sig15 vss   1.188f
C16 sig16 vss   0.208f
C25 sig25 vss   0.479f
C3  sig3  vss   0.219f
C4  sig4  vss   2.209f
C6  sig6  vss   0.436f
C12 sout  vss   0.734f
.ends
