* Tue Aug 10 11:21:07 CEST 2004
.subckt cgi2_x2 a b c vdd vss z 
*SPICE circuit <cgi2_x2> from XCircuit v3.10

m1 n4 a vss vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m2 z b n4 vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m3 n3 b vss vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m4 z c n3 vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m5 z b n2 vdd p w=74u l=2u ad='74u*5u+12p' as='74u*5u+12p' pd='74u*2+14u' ps='74u*2+14u'
m6 n2 a vdd vdd p w=74u l=2u ad='74u*5u+12p' as='74u*5u+12p' pd='74u*2+14u' ps='74u*2+14u'
m7 z c n1 vdd p w=74u l=2u ad='74u*5u+12p' as='74u*5u+12p' pd='74u*2+14u' ps='74u*2+14u'
m8 n1 b vdd vdd p w=74u l=2u ad='74u*5u+12p' as='74u*5u+12p' pd='74u*2+14u' ps='74u*2+14u'
m9 n1 a vdd vdd p w=74u l=2u ad='74u*5u+12p' as='74u*5u+12p' pd='74u*2+14u' ps='74u*2+14u'
m10 n3 a vss vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
.ends
