* Mon Aug 16 14:10:58 CEST 2004
.subckt iv1v1x2 a vdd vss z 
*SPICE circuit <iv1v1x2> from XCircuit v3.10

m1 z a vss vss n w=19u l=2.3636u ad='19u*5u+12p' as='19u*5u+12p' pd='19u*2+14u' ps='19u*2+14u'
m2 z a vdd vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
.ends
