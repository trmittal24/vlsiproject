* Spice description of rowend_x0
* Spice driver version 134999461
* Date 21/07/2007 at 19:32:27
* sxlib 0.13um values
.subckt rowend_x0 vdd vss
.ends
