magic
tech scmos
timestamp 1523032550
use empty  empty_0
timestamp 1523032550
transform 1 0 0 0 1 0
box 0 0 905 298
<< end >>
