magic
tech scmos
timestamp 1523083811
<< metal1 >>
rect 756 -387 1290 -384
rect 728 -393 1312 -390
rect 722 -401 769 -398
rect 984 -401 1030 -398
rect 1242 -400 1302 -397
rect 1309 -402 1312 -393
rect 1320 -401 1325 -398
rect 1320 -403 1324 -401
rect 1267 -411 1302 -408
rect 1245 -432 1267 -428
rect 1264 -466 1267 -432
rect 1290 -452 1293 -439
rect 1290 -456 1302 -452
rect 1264 -470 1289 -466
rect 1262 -482 1268 -478
rect 1286 -555 1289 -470
rect 1292 -548 1295 -476
rect 1292 -552 1300 -548
rect 1286 -558 1301 -555
rect 665 -587 668 -564
rect 688 -588 701 -585
rect 627 -613 631 -608
rect 698 -623 701 -588
rect 888 -612 892 -608
rect 674 -627 701 -623
rect 1195 -628 1332 -621
rect 1199 -636 1229 -633
rect 940 -656 1019 -653
rect 752 -663 763 -660
<< metal2 >>
rect 720 -378 782 -374
rect 720 -383 723 -378
rect 779 -383 782 -378
rect 970 -380 1283 -377
rect 970 -383 973 -380
rect 507 -386 723 -383
rect 507 -598 510 -386
rect 779 -386 973 -383
rect 984 -387 1276 -384
rect 752 -496 755 -387
rect 984 -396 987 -387
rect 763 -481 773 -478
rect 1023 -482 1033 -479
rect 1263 -484 1266 -411
rect 1272 -472 1276 -387
rect 1280 -443 1283 -380
rect 1290 -435 1293 -387
rect 1306 -399 1319 -397
rect 1306 -400 1316 -399
rect 1280 -447 1303 -443
rect 1272 -476 1292 -472
rect 1263 -487 1272 -484
rect 752 -499 770 -496
rect 753 -514 759 -511
rect 622 -660 625 -613
rect 622 -663 748 -660
rect 756 -669 759 -514
rect 767 -598 770 -499
rect 1269 -510 1272 -487
rect 948 -588 957 -583
rect 884 -653 887 -612
rect 884 -656 936 -653
rect 944 -660 947 -606
rect 767 -663 947 -660
rect 954 -669 957 -588
rect 756 -672 957 -669
rect 1010 -669 1013 -514
rect 1209 -588 1216 -584
rect 1027 -633 1030 -595
rect 1027 -636 1195 -633
rect 1020 -660 1023 -656
rect 1203 -660 1206 -607
rect 1020 -663 1206 -660
rect 1213 -669 1216 -588
rect 1305 -633 1308 -604
rect 1233 -636 1308 -633
rect 1010 -672 1216 -669
<< m2contact >>
rect 752 -387 756 -383
rect 1290 -387 1294 -383
rect 724 -394 728 -390
rect 1302 -400 1306 -396
rect 1316 -403 1320 -399
rect 1263 -411 1267 -407
rect 1290 -439 1294 -435
rect 759 -482 763 -478
rect 773 -482 777 -478
rect 1019 -482 1023 -478
rect 1033 -482 1037 -478
rect 749 -514 753 -510
rect 1009 -514 1013 -510
rect 1269 -514 1273 -510
rect 1292 -476 1296 -472
rect 622 -613 627 -608
rect 884 -612 888 -608
rect 1195 -636 1199 -632
rect 1229 -636 1233 -632
rect 936 -656 940 -652
rect 1019 -656 1023 -652
rect 748 -663 752 -659
rect 763 -663 767 -659
use diff2  diff2_0
timestamp 1523083811
transform 1 0 511 0 1 -473
box -4 -160 252 80
use diff2  diff2_1
timestamp 1523083811
transform 1 0 771 0 1 -473
box -4 -160 252 80
use diff2  diff2_2
timestamp 1523083811
transform 1 0 1031 0 1 -473
box -4 -160 252 80
use mux  mux_0
timestamp 1523083811
transform 1 0 1327 0 1 -473
box -29 -160 85 80
<< end >>
