* Mon Aug 16 14:22:56 CEST 2004
.subckt no2_x4 i0 i1 nq vdd vss 
*SPICE circuit <no2_x4> from XCircuit v3.10

m1 q n2 vdd vdd p w=20u l=2.3636u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m2 nq q vdd vdd p w=80u l=2.3636u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m3 n2 i1 n1 vdd p w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m4 nq q vss vss n w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m5 q n2 vss vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m6 n2 i0 vss vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m7 n2 i1 vss vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m8 n1 i0 vdd vdd p w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
.ends
