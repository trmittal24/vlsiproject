* Mon Aug 16 14:10:58 CEST 2004
.subckt iv1v0x12 a vdd vss z 
*SPICE circuit <iv1v0x12> from XCircuit v3.10

m1 z a vss vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m2 z a vdd vdd p w=160u l=2u ad='160u*5u+12p' as='160u*5u+12p' pd='160u*2+14u' ps='160u*2+14u'
.ends
