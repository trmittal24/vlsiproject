* Spice description of nr2v6x2
* Spice driver version 134999461
* Date 17/06/2007 at 14:03:27
* vgalib 0.13um values
.subckt nr2v6x2 a b vdd vss z
Mtr_00001 vss   vss   sig3  vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00002 z     a     vss   vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00003 vss   b     z     vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00004 sig5  vss   vss   vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00005 vdd   a     sig7  vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
Mtr_00006 sig7  a     vdd   vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
Mtr_00007 sig7  b     z     vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
Mtr_00008 z     b     sig7  vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
C4  a     vss   0.859f
C6  b     vss   0.870f
C7  sig7  vss   0.569f
C2  z     vss   1.024f
.ends
