* Wed Apr 11 08:42:16 CEST 2007
.subckt xor2v0x1 a b vdd vss z
*SPICE circuit <xor2v0x1> from XCircuit v3.4 rev 26

m1 z bn an vdd p w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m2 bn b vss vss n w=9u l=2u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m3 an a vss vss n w=9u l=2u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m4 n1 an vss vss n w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m5 z bn n1 vss n w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m6 an a vdd vdd p w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m7 bn b vdd vdd p w=27u l=2u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
m8 z b an vss n w=9u l=2u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m9 z an bn vdd p w=27u l=2u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
.ends
