* Thu Sep  1 18:58:46 CEST 2005
.subckt nr2v1x3 a b vdd vss z 
*SPICE circuit <nr2v1x3> from XCircuit v3.20

m1 z a vss vss n w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m2 n1 a vdd vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m3 z b vss vss n w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m4 z b n1 vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
.ends
