* Sat Mar 31 18:48:37 CEST 2007
.subckt nd2v5x3 a b vdd vss z
*SPICE circuit <nd2v5x3> from XCircuit v3.4 rev 26

m1 n1 a vss vss n w=26u l=2.3636u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m2 z a vdd vdd p w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m3 z b n1 vss n w=26u l=2.3636u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m4 z b vdd vdd p w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
.ends
