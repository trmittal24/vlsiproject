* Sat Aug 27 22:09:59 CEST 2005
.subckt iv1v4x2 a vdd vss z 
*SPICE circuit <iv1v4x2> from XCircuit v3.20

m1 z a vss vss n w=8u l=2u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
m2 z a vdd vdd p w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
.ends
