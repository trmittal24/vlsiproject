* Sun Apr  2 13:48:08 CEST 2006
.subckt or2v0x8 a b vdd vss z 
*SPICE circuit <or2v0x8> from XCircuit v3.20

m1 z zn vdd vdd p w=104u l=2.3636u ad='104u*5u+12p' as='104u*5u+12p' pd='104u*2+14u' ps='104u*2+14u'
m2 z zn vss vss n w=52u l=2.3636u ad='52u*5u+12p' as='52u*5u+12p' pd='52u*2+14u' ps='52u*2+14u'
m3 zn a vss vss n w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m4 n1 a vdd vdd p w=66u l=2.3636u ad='66u*5u+12p' as='66u*5u+12p' pd='66u*2+14u' ps='66u*2+14u'
m5 zn b vss vss n w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m6 zn b n1 vdd p w=66u l=2.3636u ad='66u*5u+12p' as='66u*5u+12p' pd='66u*2+14u' ps='66u*2+14u'
.ends
