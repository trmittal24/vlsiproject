* Tue Aug 10 11:21:07 CEST 2004
.subckt bf1_x8 a vdd vss z 
*SPICE circuit <bf1_x8> from XCircuit v3.10

m1 an a vss vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m2 an a vdd vdd p w=64u l=2u ad='64u*5u+12p' as='64u*5u+12p' pd='64u*2+14u' ps='64u*2+14u'
m3 z an vss vss n w=72u l=2u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
m4 z an vdd vdd p w=145u l=2u ad='145u*5u+12p' as='145u*5u+12p' pd='145u*2+14u' ps='145u*2+14u'
.ends
