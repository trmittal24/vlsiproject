* Spice description of vfeed5
* Spice driver version 134999461
* Date 22/07/2007 at 11:00:24
* vsxlib 0.13um values
.subckt vfeed5 vdd vss
.ends
