* Spice description of xnr2_x05
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:11
*
.subckt xnr2_x05 a b vdd vss z 
M5  vdd   a     6     vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M3  z     b     6     vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M2  n1    6     z     vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M1  vdd   sig1  n1    vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M4  sig1  b     vdd   vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M7  sig1  6     z     vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M6  z     sig1  6     vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M9  6     a     vss   vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M8  vss   b     sig1  vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
C8  a     vss   1.055f
C7  b     vss   1.115f
C6  vdd   vss   1.975f
C4  6     vss   2.875f
C3  z     vss   2.254f
C1  sig1  vss   1.572f
.ends
