* Tue Aug 10 11:21:07 CEST 2004
.subckt nr4_x1 a b c d vdd vss z 
*SPICE circuit <nr4_x1> from XCircuit v3.10

m1 z a vss vss n w=11u l=2.3636u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m2 z b vss vss n w=11u l=2.3636u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m3 z c vss vss n w=11u l=2.3636u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m4 z d vss vss n w=11u l=2.3636u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m5 z d n3 vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
m6 n3 c n2 vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
m7 n2 b n1 vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
m8 n1 a vdd vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
.ends
