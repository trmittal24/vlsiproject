magic
tech scmos
timestamp 1523084160
use totdiff3  totdiff3_0
timestamp 1523084160
transform 1 0 -569 0 1 937
box 507 -672 1412 -374
use ../../../../prac/counter  counter_0 ../../../../prac
timestamp 1523084160
transform 1 0 608 0 1 76
box -608 -76 216 157
<< end >>
