* SPICE3 file created from final.ext - technology: scmos

.option scale=1u

M1000 3seg_0/2seg_0/an2v0x3_0/a 3seg_0/2seg_0/or3v0x3_0/zn vdd vdd pfet w=19 l=2
+ ad=162 pd=58 as=35339 ps=12852 
M1001 vdd 3seg_0/2seg_0/or3v0x3_0/zn 3seg_0/2seg_0/an2v0x3_0/a vdd pfet w=21 l=2
+ ad=0 pd=0 as=0 ps=0 
M1002 3seg_0/2seg_0/or3v0x3_0/a_33_38# 3seg_0/2seg_0/or3v0x3_0/a vdd vdd pfet w=28 l=2
+ ad=140 pd=66 as=0 ps=0 
M1003 3seg_0/2seg_0/or3v0x3_0/a_40_38# 3seg_0/2seg_0/or3v0x3_0/b 3seg_0/2seg_0/or3v0x3_0/a_33_38# vdd pfet w=28 l=2
+ ad=140 pd=66 as=0 ps=0 
M1004 3seg_0/2seg_0/or3v0x3_0/zn 3seg_0/2seg_0/or3v0x3_0/c 3seg_0/2seg_0/or3v0x3_0/a_40_38# vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1005 3seg_0/2seg_0/or3v0x3_0/a_57_38# 3seg_0/2seg_0/or3v0x3_0/c 3seg_0/2seg_0/or3v0x3_0/zn vdd pfet w=28 l=2
+ ad=140 pd=66 as=0 ps=0 
M1006 3seg_0/2seg_0/or3v0x3_0/a_64_38# 3seg_0/2seg_0/or3v0x3_0/b 3seg_0/2seg_0/or3v0x3_0/a_57_38# vdd pfet w=28 l=2
+ ad=140 pd=66 as=0 ps=0 
M1007 vdd 3seg_0/2seg_0/or3v0x3_0/a 3seg_0/2seg_0/or3v0x3_0/a_64_38# vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1008 gnd 3seg_0/2seg_0/or3v0x3_0/zn 3seg_0/2seg_0/an2v0x3_0/a gnd nfet w=20 l=2
+ ad=25596 pd=8510 as=126 ps=54 
M1009 3seg_0/2seg_0/or3v0x3_0/zn 3seg_0/2seg_0/or3v0x3_0/a gnd gnd nfet w=10 l=2
+ ad=142 pd=70 as=0 ps=0 
M1010 gnd 3seg_0/2seg_0/or3v0x3_0/b 3seg_0/2seg_0/or3v0x3_0/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1011 3seg_0/2seg_0/or3v0x3_0/zn 3seg_0/2seg_0/or3v0x3_0/c gnd gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1012 3seg_0/2seg_0/an2v0x3_0/z 3seg_0/2seg_0/an2v0x3_0/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1013 vdd 3seg_0/2seg_0/an2v0x3_0/zn 3seg_0/2seg_0/an2v0x3_0/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1014 3seg_0/2seg_0/an2v0x3_0/zn 3seg_0/2seg_0/an2v0x3_0/a vdd vdd pfet w=20 l=2
+ ad=166 pd=62 as=0 ps=0 
M1015 vdd 3seg_0/2seg_0/an2v0x3_0/b 3seg_0/2seg_0/an2v0x3_0/zn vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1016 gnd 3seg_0/2seg_0/an2v0x3_0/zn 3seg_0/2seg_0/an2v0x3_0/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1017 3seg_0/2seg_0/an2v0x3_0/a_30_9# 3seg_0/2seg_0/an2v0x3_0/a gnd gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1018 3seg_0/2seg_0/an2v0x3_0/zn 3seg_0/2seg_0/an2v0x3_0/b 3seg_0/2seg_0/an2v0x3_0/a_30_9# gnd nfet w=17 l=2
+ ad=97 pd=48 as=0 ps=0 
M1019 3seg_0/2seg_0/1counter_0/an2v0x3_1/b 3seg_0/2seg_0/ud vdd vdd pfet w=24 l=2
+ ad=168 pd=64 as=0 ps=0 
M1020 vdd 3seg_0/2seg_0/ud 3seg_0/2seg_0/1counter_0/an2v0x3_1/b vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1021 3seg_0/2seg_0/1counter_0/an2v0x3_1/b 3seg_0/2seg_0/ud gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1022 gnd 3seg_0/2seg_0/ud 3seg_0/2seg_0/1counter_0/an2v0x3_1/b gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1023 3seg_0/2seg_0/1counter_0/an2v0x3_2/b 3seg_0/2seg_0/1counter_0/an2v0x3_1/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1024 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_1/zn 3seg_0/2seg_0/1counter_0/an2v0x3_2/b vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1025 3seg_0/2seg_0/1counter_0/an2v0x3_1/zn 3seg_0/2seg_0/1counter_0/an2v0x3_1/a vdd vdd pfet w=20 l=2
+ ad=166 pd=62 as=0 ps=0 
M1026 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_1/b 3seg_0/2seg_0/1counter_0/an2v0x3_1/zn vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1027 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_1/zn 3seg_0/2seg_0/1counter_0/an2v0x3_2/b gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1028 3seg_0/2seg_0/1counter_0/an2v0x3_1/a_30_9# 3seg_0/2seg_0/1counter_0/an2v0x3_1/a gnd gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1029 3seg_0/2seg_0/1counter_0/an2v0x3_1/zn 3seg_0/2seg_0/1counter_0/an2v0x3_1/b 3seg_0/2seg_0/1counter_0/an2v0x3_1/a_30_9# gnd nfet w=17 l=2
+ ad=97 pd=48 as=0 ps=0 
M1030 3seg_0/2seg_0/1counter_0/an2v0x3_2/z 3seg_0/2seg_0/1counter_0/an2v0x3_2/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1031 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_2/zn 3seg_0/2seg_0/1counter_0/an2v0x3_2/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1032 3seg_0/2seg_0/1counter_0/an2v0x3_2/zn 3seg_0/2seg_0/1counter_0/an2v0x3_2/a vdd vdd pfet w=20 l=2
+ ad=166 pd=62 as=0 ps=0 
M1033 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_2/b 3seg_0/2seg_0/1counter_0/an2v0x3_2/zn vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1034 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_2/zn 3seg_0/2seg_0/1counter_0/an2v0x3_2/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1035 3seg_0/2seg_0/1counter_0/an2v0x3_2/a_30_9# 3seg_0/2seg_0/1counter_0/an2v0x3_2/a gnd gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1036 3seg_0/2seg_0/1counter_0/an2v0x3_2/zn 3seg_0/2seg_0/1counter_0/an2v0x3_2/b 3seg_0/2seg_0/1counter_0/an2v0x3_2/a_30_9# gnd nfet w=17 l=2
+ ad=97 pd=48 as=0 ps=0 
M1037 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/a 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/bn vdd pfet w=21 l=2
+ ad=0 pd=0 as=248 ps=112 
M1038 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/an 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/a vdd vdd pfet w=13 l=2
+ ad=104 pd=42 as=0 ps=0 
M1039 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/bn 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/an vdd pfet w=13 l=2
+ ad=144 pd=58 as=0 ps=0 
M1040 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/bn 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/an 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/d vdd pfet w=21 l=2
+ ad=0 pd=0 as=0 ps=0 
M1041 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/a 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/bn gnd nfet w=7 l=2
+ ad=0 pd=0 as=49 ps=28 
M1042 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/an 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/a gnd gnd nfet w=7 l=2
+ ad=56 pd=30 as=0 ps=0 
M1043 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/bf1v0x4_0/a 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/an gnd nfet w=7 l=2
+ ad=66 pd=34 as=0 ps=0 
M1044 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/a_48_11# 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/bn 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/d gnd nfet w=9 l=2
+ ad=45 pd=28 as=0 ps=0 
M1045 gnd 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/an 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/a_48_11# gnd nfet w=9 l=2
+ ad=0 pd=0 as=0 ps=0 
M1046 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_1/a 3seg_0/2seg_0/1counter_0/bf1v0x4_0/a vdd pfet w=28 l=2
+ ad=0 pd=0 as=168 ps=70 
M1047 3seg_0/2seg_0/1counter_0/an2v0x3_1/a 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n4 vdd vdd pfet w=14 l=2
+ ad=82 pd=42 as=0 ps=0 
M1048 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/a_40_48# 3seg_0/2seg_0/1counter_0/an2v0x3_1/a vdd vdd pfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1049 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n4 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/a_40_48# vdd pfet w=6 l=2
+ ad=78 pd=40 as=0 ps=0 
M1050 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n2 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n4 vdd pfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1051 vdd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n1 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n2 vdd pfet w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1052 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/a_77_54# 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n2 vdd vdd pfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1053 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n1 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/a_77_54# vdd pfet w=6 l=2
+ ad=83 pd=42 as=0 ps=0 
M1054 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_1/a 3seg_0/2seg_0/1counter_0/bf1v0x4_0/a gnd nfet w=14 l=2
+ ad=0 pd=0 as=82 ps=42 
M1055 gnd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n4 3seg_0/2seg_0/1counter_0/an2v0x3_1/a gnd nfet w=7 l=2
+ ad=0 pd=0 as=47 ps=28 
M1056 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/a_94_47# 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n1 vdd pfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1057 vdd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/a_94_47# vdd pfet w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1058 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/cn vdd vdd pfet w=11 l=2
+ ad=67 pd=36 as=0 ps=0 
M1059 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/cn 3seg_0/2seg_0/an2v0x3_0/z vdd vdd pfet w=10 l=2
+ ad=62 pd=34 as=0 ps=0 
M1060 gnd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/ci gnd nfet w=6 l=2
+ ad=0 pd=0 as=42 ps=26 
M1061 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/a_40_13# 3seg_0/2seg_0/1counter_0/an2v0x3_1/a gnd gnd nfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1062 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n4 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/a_40_13# gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1063 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n2 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n4 gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1064 gnd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n1 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n2 gnd nfet w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1065 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/a_77_13# 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n2 gnd gnd nfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1066 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n1 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/a_77_13# gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1067 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/a_94_13# 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n1 gnd nfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1068 gnd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/a_94_13# gnd nfet w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1069 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/cn 3seg_0/2seg_0/an2v0x3_0/z gnd gnd nfet w=7 l=2
+ ad=49 pd=28 as=0 ps=0 
M1070 3seg_0/2seg_0/1counter_0/or2v0x3_0/z 3seg_0/2seg_0/1counter_0/or2v0x3_0/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1071 vdd 3seg_0/2seg_0/1counter_0/or2v0x3_0/zn 3seg_0/2seg_0/1counter_0/or2v0x3_0/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1072 3seg_0/2seg_0/1counter_0/or2v0x3_0/a_31_39# 3seg_0/2seg_0/1counter_0/an2v0x3_3/b vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1073 3seg_0/2seg_0/1counter_0/or2v0x3_0/zn 3seg_0/2seg_0/1counter_0/an2v0x3_2/b 3seg_0/2seg_0/1counter_0/or2v0x3_0/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1074 3seg_0/2seg_0/1counter_0/or2v0x3_0/a_48_39# 3seg_0/2seg_0/1counter_0/an2v0x3_2/b 3seg_0/2seg_0/1counter_0/or2v0x3_0/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1075 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_3/b 3seg_0/2seg_0/1counter_0/or2v0x3_0/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1076 gnd 3seg_0/2seg_0/1counter_0/or2v0x3_0/zn 3seg_0/2seg_0/1counter_0/or2v0x3_0/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1077 3seg_0/2seg_0/1counter_0/or2v0x3_0/zn 3seg_0/2seg_0/1counter_0/an2v0x3_3/b gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1078 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_2/b 3seg_0/2seg_0/1counter_0/or2v0x3_0/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1079 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/bn vdd pfet w=21 l=2
+ ad=0 pd=0 as=248 ps=112 
M1080 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/an 3seg_0/2seg_0/1counter_0/or2v0x3_0/z vdd vdd pfet w=13 l=2
+ ad=104 pd=42 as=0 ps=0 
M1081 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/bn 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/an vdd pfet w=13 l=2
+ ad=144 pd=58 as=0 ps=0 
M1082 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/bn 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/an 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/d vdd pfet w=21 l=2
+ ad=0 pd=0 as=0 ps=0 
M1083 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/bn gnd nfet w=7 l=2
+ ad=0 pd=0 as=49 ps=28 
M1084 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/an 3seg_0/2seg_0/1counter_0/or2v0x3_0/z gnd gnd nfet w=7 l=2
+ ad=56 pd=30 as=0 ps=0 
M1085 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/an gnd nfet w=7 l=2
+ ad=66 pd=34 as=0 ps=0 
M1086 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/a_48_11# 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/bn 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/d gnd nfet w=9 l=2
+ ad=45 pd=28 as=0 ps=0 
M1087 gnd 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/an 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/a_48_11# gnd nfet w=9 l=2
+ ad=0 pd=0 as=0 ps=0 
M1088 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_2/a 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a vdd pfet w=28 l=2
+ ad=0 pd=0 as=168 ps=70 
M1089 3seg_0/2seg_0/1counter_0/an2v0x3_2/a 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n4 vdd vdd pfet w=14 l=2
+ ad=82 pd=42 as=0 ps=0 
M1090 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/a_40_48# 3seg_0/2seg_0/1counter_0/an2v0x3_2/a vdd vdd pfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1091 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n4 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/a_40_48# vdd pfet w=6 l=2
+ ad=78 pd=40 as=0 ps=0 
M1092 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n2 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n4 vdd pfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1093 vdd 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n1 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n2 vdd pfet w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1094 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/a_77_54# 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n2 vdd vdd pfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1095 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n1 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/a_77_54# vdd pfet w=6 l=2
+ ad=83 pd=42 as=0 ps=0 
M1096 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_2/a 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a gnd nfet w=14 l=2
+ ad=0 pd=0 as=82 ps=42 
M1097 gnd 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n4 3seg_0/2seg_0/1counter_0/an2v0x3_2/a gnd nfet w=7 l=2
+ ad=0 pd=0 as=47 ps=28 
M1098 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/a_94_47# 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n1 vdd pfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1099 vdd 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/a_94_47# vdd pfet w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1100 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/cn vdd vdd pfet w=11 l=2
+ ad=67 pd=36 as=0 ps=0 
M1101 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/cn 3seg_0/2seg_0/an2v0x3_0/z vdd vdd pfet w=10 l=2
+ ad=62 pd=34 as=0 ps=0 
M1102 gnd 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/ci gnd nfet w=6 l=2
+ ad=0 pd=0 as=42 ps=26 
M1103 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/a_40_13# 3seg_0/2seg_0/1counter_0/an2v0x3_2/a gnd gnd nfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1104 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n4 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/a_40_13# gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1105 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n2 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n4 gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1106 gnd 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n1 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n2 gnd nfet w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1107 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/a_77_13# 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n2 gnd gnd nfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1108 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n1 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/a_77_13# gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1109 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/a_94_13# 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n1 gnd nfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1110 gnd 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/a_94_13# gnd nfet w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1111 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/cn 3seg_0/2seg_0/an2v0x3_0/z gnd gnd nfet w=7 l=2
+ ad=49 pd=28 as=0 ps=0 
M1112 3seg_0/2seg_0/1counter_0/or2v0x3_1/z 3seg_0/2seg_0/1counter_0/or2v0x3_1/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1113 vdd 3seg_0/2seg_0/1counter_0/or2v0x3_1/zn 3seg_0/2seg_0/1counter_0/or2v0x3_1/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1114 3seg_0/2seg_0/1counter_0/or2v0x3_1/a_31_39# 3seg_0/2seg_0/1counter_0/or2v0x3_1/a vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1115 3seg_0/2seg_0/1counter_0/or2v0x3_1/zn 3seg_0/2seg_0/1counter_0/an2v0x3_2/z 3seg_0/2seg_0/1counter_0/or2v0x3_1/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1116 3seg_0/2seg_0/1counter_0/or2v0x3_1/a_48_39# 3seg_0/2seg_0/1counter_0/an2v0x3_2/z 3seg_0/2seg_0/1counter_0/or2v0x3_1/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1117 vdd 3seg_0/2seg_0/1counter_0/or2v0x3_1/a 3seg_0/2seg_0/1counter_0/or2v0x3_1/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1118 gnd 3seg_0/2seg_0/1counter_0/or2v0x3_1/zn 3seg_0/2seg_0/1counter_0/or2v0x3_1/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1119 3seg_0/2seg_0/1counter_0/or2v0x3_1/zn 3seg_0/2seg_0/1counter_0/or2v0x3_1/a gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1120 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_2/z 3seg_0/2seg_0/1counter_0/or2v0x3_1/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1121 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/a 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/bn vdd pfet w=21 l=2
+ ad=0 pd=0 as=248 ps=112 
M1122 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/an 3seg_0/2seg_0/1counter_0/or2v0x3_1/z vdd vdd pfet w=13 l=2
+ ad=104 pd=42 as=0 ps=0 
M1123 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/bn 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/an vdd pfet w=13 l=2
+ ad=144 pd=58 as=0 ps=0 
M1124 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/bn 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/an 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/d vdd pfet w=21 l=2
+ ad=0 pd=0 as=0 ps=0 
M1125 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/a 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/bn gnd nfet w=7 l=2
+ ad=0 pd=0 as=49 ps=28 
M1126 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/an 3seg_0/2seg_0/1counter_0/or2v0x3_1/z gnd gnd nfet w=7 l=2
+ ad=56 pd=30 as=0 ps=0 
M1127 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/bf1v0x4_2/a 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/an gnd nfet w=7 l=2
+ ad=66 pd=34 as=0 ps=0 
M1128 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/a_48_11# 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/bn 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/d gnd nfet w=9 l=2
+ ad=45 pd=28 as=0 ps=0 
M1129 gnd 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/an 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/a_48_11# gnd nfet w=9 l=2
+ ad=0 pd=0 as=0 ps=0 
M1130 vdd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/zn 3seg_0/2seg_0/1counter_0/bf1v0x4_2/a vdd pfet w=28 l=2
+ ad=0 pd=0 as=168 ps=70 
M1131 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/zn 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n4 vdd vdd pfet w=14 l=2
+ ad=82 pd=42 as=0 ps=0 
M1132 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/a_40_48# 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/zn vdd vdd pfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1133 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n4 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/a_40_48# vdd pfet w=6 l=2
+ ad=78 pd=40 as=0 ps=0 
M1134 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n2 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n4 vdd pfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1135 vdd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n1 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n2 vdd pfet w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1136 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/a_77_54# 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n2 vdd vdd pfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1137 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n1 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/a_77_54# vdd pfet w=6 l=2
+ ad=83 pd=42 as=0 ps=0 
M1138 gnd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/zn 3seg_0/2seg_0/1counter_0/bf1v0x4_2/a gnd nfet w=14 l=2
+ ad=0 pd=0 as=82 ps=42 
M1139 gnd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n4 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/zn gnd nfet w=7 l=2
+ ad=0 pd=0 as=47 ps=28 
M1140 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/a_94_47# 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n1 vdd pfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1141 vdd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/a_94_47# vdd pfet w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1142 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/cn vdd vdd pfet w=11 l=2
+ ad=67 pd=36 as=0 ps=0 
M1143 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/cn 3seg_0/2seg_0/an2v0x3_0/z vdd vdd pfet w=10 l=2
+ ad=62 pd=34 as=0 ps=0 
M1144 gnd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/ci gnd nfet w=6 l=2
+ ad=0 pd=0 as=42 ps=26 
M1145 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/a_40_13# 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/zn gnd gnd nfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1146 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n4 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/a_40_13# gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1147 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n2 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n4 gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1148 gnd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n1 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n2 gnd nfet w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1149 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/a_77_13# 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n2 gnd gnd nfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1150 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n1 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/a_77_13# gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1151 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/a_94_13# 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/cn 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n1 gnd nfet w=6 l=2
+ ad=30 pd=22 as=0 ps=0 
M1152 gnd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/a_94_13# gnd nfet w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1153 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/cn 3seg_0/2seg_0/an2v0x3_0/z gnd gnd nfet w=7 l=2
+ ad=49 pd=28 as=0 ps=0 
M1154 3seg_0/2seg_0/1counter_0/an2v0x3_3/b 3seg_0/2seg_0/1counter_0/an2v0x3_0/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1155 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_0/zn 3seg_0/2seg_0/1counter_0/an2v0x3_3/b vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1156 3seg_0/2seg_0/1counter_0/an2v0x3_0/zn 3seg_0/2seg_0/ud vdd vdd pfet w=20 l=2
+ ad=166 pd=62 as=0 ps=0 
M1157 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z 3seg_0/2seg_0/1counter_0/an2v0x3_0/zn vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1158 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_0/zn 3seg_0/2seg_0/1counter_0/an2v0x3_3/b gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1159 3seg_0/2seg_0/1counter_0/an2v0x3_0/a_30_9# 3seg_0/2seg_0/ud gnd gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1160 3seg_0/2seg_0/1counter_0/an2v0x3_0/zn 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z 3seg_0/2seg_0/1counter_0/an2v0x3_0/a_30_9# gnd nfet w=17 l=2
+ ad=97 pd=48 as=0 ps=0 
M1161 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z 3seg_0/2seg_0/1counter_0/bf1v0x4_0/an vdd vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1162 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/an 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1163 3seg_0/2seg_0/1counter_0/bf1v0x4_0/an 3seg_0/2seg_0/1counter_0/bf1v0x4_0/a vdd vdd pfet w=27 l=2
+ ad=161 pd=68 as=0 ps=0 
M1164 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z 3seg_0/2seg_0/1counter_0/bf1v0x4_0/an gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/w_n4_n4# nfet w=14 l=2
+ ad=112 pd=44 as=0 ps=0 
M1165 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/an 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z 3seg_0/2seg_0/1counter_0/bf1v0x4_0/w_n4_n4# nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1166 3seg_0/2seg_0/1counter_0/bf1v0x4_0/an 3seg_0/2seg_0/1counter_0/bf1v0x4_0/a gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/w_n4_n4# nfet w=15 l=2
+ ad=101 pd=44 as=0 ps=0 
M1167 3seg_0/2seg_0/1counter_0/or2v0x3_1/a 3seg_0/2seg_0/1counter_0/an2v0x3_3/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1168 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_3/zn 3seg_0/2seg_0/1counter_0/or2v0x3_1/a vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1169 3seg_0/2seg_0/1counter_0/an2v0x3_3/zn 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z vdd vdd pfet w=20 l=2
+ ad=166 pd=62 as=0 ps=0 
M1170 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_3/b 3seg_0/2seg_0/1counter_0/an2v0x3_3/zn vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1171 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_3/zn 3seg_0/2seg_0/1counter_0/or2v0x3_1/a gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1172 3seg_0/2seg_0/1counter_0/an2v0x3_3/a_30_9# 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z gnd gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1173 3seg_0/2seg_0/1counter_0/an2v0x3_3/zn 3seg_0/2seg_0/1counter_0/an2v0x3_3/b 3seg_0/2seg_0/1counter_0/an2v0x3_3/a_30_9# gnd nfet w=17 l=2
+ ad=97 pd=48 as=0 ps=0 
M1174 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z 3seg_0/2seg_0/1counter_0/bf1v0x4_1/an vdd vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1175 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_1/an 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1176 3seg_0/2seg_0/1counter_0/bf1v0x4_1/an 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a vdd vdd pfet w=27 l=2
+ ad=161 pd=68 as=0 ps=0 
M1177 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z 3seg_0/2seg_0/1counter_0/bf1v0x4_1/an gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_1/w_n4_n4# nfet w=14 l=2
+ ad=112 pd=44 as=0 ps=0 
M1178 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_1/an 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z 3seg_0/2seg_0/1counter_0/bf1v0x4_1/w_n4_n4# nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1179 3seg_0/2seg_0/1counter_0/bf1v0x4_1/an 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_1/w_n4_n4# nfet w=15 l=2
+ ad=101 pd=44 as=0 ps=0 
M1180 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z 3seg_0/2seg_0/1counter_0/bf1v0x4_2/an vdd vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1181 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/an 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1182 3seg_0/2seg_0/1counter_0/bf1v0x4_2/an 3seg_0/2seg_0/1counter_0/bf1v0x4_2/a vdd vdd pfet w=27 l=2
+ ad=161 pd=68 as=0 ps=0 
M1183 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z 3seg_0/2seg_0/1counter_0/bf1v0x4_2/an gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/w_n4_n4# nfet w=14 l=2
+ ad=112 pd=44 as=0 ps=0 
M1184 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/an 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z 3seg_0/2seg_0/1counter_0/bf1v0x4_2/w_n4_n4# nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1185 3seg_0/2seg_0/1counter_0/bf1v0x4_2/an 3seg_0/2seg_0/1counter_0/bf1v0x4_2/a gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/w_n4_n4# nfet w=15 l=2
+ ad=101 pd=44 as=0 ps=0 
M1186 3seg_0/2seg_0/iv1v0x3_0/z 3seg_0/2seg_0/iv1v0x3_0/a vdd vdd pfet w=24 l=2
+ ad=168 pd=64 as=0 ps=0 
M1187 vdd 3seg_0/2seg_0/iv1v0x3_0/a 3seg_0/2seg_0/iv1v0x3_0/z vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1188 3seg_0/2seg_0/iv1v0x3_0/z 3seg_0/2seg_0/iv1v0x3_0/a gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1189 gnd 3seg_0/2seg_0/iv1v0x3_0/a 3seg_0/2seg_0/iv1v0x3_0/z gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1190 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/zn 3seg_0/2seg_0/or3v0x3_0/c 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# pfet w=18 l=2
+ ad=0 pd=0 as=102 ps=50 
M1191 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/a_21_50# 3seg_0/2seg_0/totdiff3_0/mux_0/a2 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1192 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/zn 3seg_0/2seg_0/ud 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/a_21_50# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=128 pd=48 as=0 ps=0 
M1193 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/a_38_50# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/sn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/zn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1194 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/b2 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/a_38_50# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1195 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/sn 3seg_0/2seg_0/ud vdd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# pfet w=8 l=2
+ ad=52 pd=30 as=0 ps=0 
M1196 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/zn 3seg_0/2seg_0/or3v0x3_0/c 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# nfet w=9 l=2
+ ad=0 pd=0 as=57 ps=32 
M1197 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/a_21_12# 3seg_0/2seg_0/totdiff3_0/mux_0/a2 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# nfet w=8 l=2
+ ad=40 pd=26 as=0 ps=0 
M1198 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/zn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/sn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/a_21_12# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# nfet w=8 l=2
+ ad=64 pd=32 as=0 ps=0 
M1199 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/a_38_12# 3seg_0/2seg_0/ud 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/zn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# nfet w=8 l=2
+ ad=40 pd=26 as=0 ps=0 
M1200 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/b2 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/a_38_12# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1201 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/sn 3seg_0/2seg_0/ud gnd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# nfet w=6 l=2
+ ad=42 pd=26 as=0 ps=0 
M1202 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/zn 3seg_0/2seg_0/or3v0x3_0/b 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# pfet w=18 l=2
+ ad=0 pd=0 as=102 ps=50 
M1203 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/a_21_50# 3seg_0/2seg_0/totdiff3_0/mux_0/a1 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1204 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/zn 3seg_0/2seg_0/ud 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/a_21_50# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=128 pd=48 as=0 ps=0 
M1205 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/a_38_50# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/sn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/zn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1206 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/b1 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/a_38_50# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1207 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/sn 3seg_0/2seg_0/ud vdd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# pfet w=8 l=2
+ ad=52 pd=30 as=0 ps=0 
M1208 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/zn 3seg_0/2seg_0/or3v0x3_0/b 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# nfet w=9 l=2
+ ad=0 pd=0 as=57 ps=32 
M1209 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/a_21_12# 3seg_0/2seg_0/totdiff3_0/mux_0/a1 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=40 pd=26 as=0 ps=0 
M1210 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/zn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/sn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/a_21_12# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=64 pd=32 as=0 ps=0 
M1211 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/a_38_12# 3seg_0/2seg_0/ud 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/zn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=40 pd=26 as=0 ps=0 
M1212 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/b1 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/a_38_12# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1213 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/sn 3seg_0/2seg_0/ud gnd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# nfet w=6 l=2
+ ad=42 pd=26 as=0 ps=0 
M1214 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/zn 3seg_0/2seg_0/or3v0x3_0/a 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# pfet w=18 l=2
+ ad=0 pd=0 as=102 ps=50 
M1215 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/a_21_50# 3seg_0/2seg_0/totdiff3_0/mux_0/a0 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1216 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/zn 3seg_0/2seg_0/ud 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/a_21_50# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# pfet w=16 l=2
+ ad=128 pd=48 as=0 ps=0 
M1217 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/a_38_50# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/sn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/zn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1218 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/b0 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/a_38_50# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1219 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/sn 3seg_0/2seg_0/ud vdd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# pfet w=8 l=2
+ ad=52 pd=30 as=0 ps=0 
M1220 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/zn 3seg_0/2seg_0/or3v0x3_0/a 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# nfet w=9 l=2
+ ad=0 pd=0 as=57 ps=32 
M1221 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/a_21_12# 3seg_0/2seg_0/totdiff3_0/mux_0/a0 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=40 pd=26 as=0 ps=0 
M1222 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/zn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/sn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/a_21_12# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=64 pd=32 as=0 ps=0 
M1223 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/a_38_12# 3seg_0/2seg_0/ud 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/zn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=40 pd=26 as=0 ps=0 
M1224 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/b0 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/a_38_12# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1225 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/sn 3seg_0/2seg_0/ud gnd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# nfet w=6 l=2
+ ad=42 pd=26 as=0 ps=0 
M1226 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1227 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1228 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/in_2c 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1229 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1230 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a_24_13# 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1231 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/in_2c 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1232 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/mux_0/b2 vdd pfet w=20 l=2
+ ad=320 pd=112 as=398 ps=164 
M1233 3seg_0/2seg_0/totdiff3_0/mux_0/b2 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1234 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/mux_0/b2 vdd pfet w=20 l=2
+ ad=320 pd=112 as=0 ps=0 
M1235 3seg_0/2seg_0/totdiff3_0/mux_0/b2 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1236 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_2/in_2c vdd vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1237 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/in_2c 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1238 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a vdd vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1239 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1240 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/a_13_13# 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1241 3seg_0/2seg_0/totdiff3_0/mux_0/b2 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/a_13_13# gnd nfet w=13 l=2
+ ad=264 pd=98 as=0 ps=0 
M1242 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/a_30_13# 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/mux_0/b2 gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1243 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/a_30_13# gnd nfet w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1244 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_2/in_2c gnd gnd nfet w=10 l=2
+ ad=130 pd=56 as=0 ps=0 
M1245 3seg_0/2seg_0/totdiff3_0/mux_0/b2 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn gnd nfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1246 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_2/in_2c 3seg_0/2seg_0/totdiff3_0/mux_0/b2 gnd nfet w=20 l=2
+ ad=130 pd=56 as=0 ps=0 
M1247 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1248 3seg_0/2seg_0/ud 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1249 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/zn 3seg_0/2seg_0/ud vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1250 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/a_31_39# 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/z vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1251 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/z 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1252 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/a_48_39# 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/z 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1253 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/z 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1254 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/zn 3seg_0/2seg_0/ud gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1255 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/z gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1256 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/z 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1257 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1258 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1259 vdd 3seg_0/firseg_0/3_bitmux_0/o2 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1260 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1261 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a_24_13# 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1262 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/zn 3seg_0/firseg_0/3_bitmux_0/o2 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1263 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1264 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1265 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/b 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1266 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1267 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/a_24_13# 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1268 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/b 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1269 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/b vdd pfet w=12 l=2
+ ad=0 pd=0 as=72 ps=38 
M1270 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/an 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z vdd vdd pfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1271 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/an vdd pfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1272 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/ai 3seg_0/firseg_0/3_bitmux_0/o2 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/zn vdd pfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1273 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/an 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/ai vdd pfet w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1274 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/bn 3seg_0/firseg_0/3_bitmux_0/o2 vdd vdd pfet w=12 l=2
+ ad=72 pd=38 as=0 ps=0 
M1275 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/b gnd nfet w=6 l=2
+ ad=0 pd=0 as=42 ps=26 
M1276 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/an 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z gnd gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1277 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/zn 3seg_0/firseg_0/3_bitmux_0/o2 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/an gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1278 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/ai 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/zn gnd nfet w=6 l=2
+ ad=57 pd=32 as=0 ps=0 
M1279 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/an 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/ai gnd nfet w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1280 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/bn 3seg_0/firseg_0/3_bitmux_0/o2 gnd gnd nfet w=6 l=2
+ ad=42 pd=26 as=0 ps=0 
M1281 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/mux_0/a2 vdd vdd pfet w=24 l=2
+ ad=168 pd=64 as=0 ps=0 
M1282 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/a2 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1283 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/mux_0/a2 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1284 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/a2 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1285 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/mux_0/a2 vdd pfet w=27 l=2
+ ad=424 pd=138 as=530 ps=208 
M1286 3seg_0/2seg_0/totdiff3_0/mux_0/a2 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn vdd pfet w=27 l=2
+ ad=0 pd=0 as=0 ps=0 
M1287 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/mux_0/a2 vdd pfet w=27 l=2
+ ad=440 pd=142 as=0 ps=0 
M1288 3seg_0/2seg_0/totdiff3_0/mux_0/a2 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn vdd pfet w=27 l=2
+ ad=0 pd=0 as=0 ps=0 
M1289 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c vdd vdd pfet w=26 l=2
+ ad=0 pd=0 as=0 ps=0 
M1290 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn vdd pfet w=26 l=2
+ ad=0 pd=0 as=0 ps=0 
M1291 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/iz vdd vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1292 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1293 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/bn vdd pfet w=28 l=2
+ ad=224 pd=72 as=272 ps=122 
M1294 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/iz vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1295 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1296 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/bn 3seg_0/firseg_0/3_bitmux_0/o2 vdd vdd pfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1297 vdd 3seg_0/firseg_0/3_bitmux_0/o2 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/bn vdd pfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1298 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/a_11_12# 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn gnd gnd nfet w=12 l=2
+ ad=60 pd=34 as=0 ps=0 
M1299 3seg_0/2seg_0/totdiff3_0/mux_0/a2 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/a_11_12# gnd nfet w=12 l=2
+ ad=208 pd=84 as=0 ps=0 
M1300 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/a_28_12# 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/mux_0/a2 gnd nfet w=12 l=2
+ ad=60 pd=34 as=0 ps=0 
M1301 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/a_28_12# gnd nfet w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1302 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/iz gnd gnd nfet w=14 l=2
+ ad=224 pd=88 as=0 ps=0 
M1303 3seg_0/2seg_0/totdiff3_0/mux_0/a2 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn gnd nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1304 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c 3seg_0/2seg_0/totdiff3_0/mux_0/a2 gnd nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1305 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn gnd nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1306 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c gnd gnd nfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1307 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn gnd nfet w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1308 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/a_115_7# 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1309 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/a_115_7# gnd nfet w=13 l=2
+ ad=104 pd=42 as=0 ps=0 
M1310 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a 3seg_0/firseg_0/3_bitmux_0/o2 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/iz gnd nfet w=13 l=2
+ ad=114 pd=52 as=0 ps=0 
M1311 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a gnd nfet w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1312 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/bn 3seg_0/firseg_0/3_bitmux_0/o2 gnd gnd nfet w=11 l=2
+ ad=67 pd=36 as=0 ps=0 
M1313 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/in_2c vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1314 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1315 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/in_2c 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1316 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/in_2c gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1317 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a_24_13# 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1318 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/in_2c 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1319 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/mux_0/b1 vdd pfet w=20 l=2
+ ad=320 pd=112 as=398 ps=164 
M1320 3seg_0/2seg_0/totdiff3_0/mux_0/b1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1321 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/mux_0/b1 vdd pfet w=20 l=2
+ ad=320 pd=112 as=0 ps=0 
M1322 3seg_0/2seg_0/totdiff3_0/mux_0/b1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1323 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_1/in_2c vdd vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1324 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/in_2c 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1325 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a vdd vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1326 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1327 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/a_13_13# 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1328 3seg_0/2seg_0/totdiff3_0/mux_0/b1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/a_13_13# gnd nfet w=13 l=2
+ ad=264 pd=98 as=0 ps=0 
M1329 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/a_30_13# 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/mux_0/b1 gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1330 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/a_30_13# gnd nfet w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1331 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_1/in_2c gnd gnd nfet w=10 l=2
+ ad=130 pd=56 as=0 ps=0 
M1332 3seg_0/2seg_0/totdiff3_0/mux_0/b1 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn gnd nfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1333 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_1/in_2c 3seg_0/2seg_0/totdiff3_0/mux_0/b1 gnd nfet w=20 l=2
+ ad=130 pd=56 as=0 ps=0 
M1334 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1335 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1336 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1337 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/a_31_39# 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/z vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1338 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/z 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1339 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/a_48_39# 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/z 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1340 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/z 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1341 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1342 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/z gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1343 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/z 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1344 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1345 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1346 vdd 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1347 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1348 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a_24_13# 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1349 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/zn 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1350 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1351 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1352 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/b 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1353 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1354 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/a_24_13# 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1355 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/b 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1356 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/b vdd pfet w=12 l=2
+ ad=0 pd=0 as=72 ps=38 
M1357 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/an 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z vdd vdd pfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1358 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/an vdd pfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1359 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/ai 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/zn vdd pfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1360 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/an 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/ai vdd pfet w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1361 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/bn 3seg_0/firseg_0/3_bitmux_0/o1 vdd vdd pfet w=12 l=2
+ ad=72 pd=38 as=0 ps=0 
M1362 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/b gnd nfet w=6 l=2
+ ad=0 pd=0 as=42 ps=26 
M1363 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/an 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z gnd gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1364 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/zn 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/an gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1365 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/ai 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/zn gnd nfet w=6 l=2
+ ad=57 pd=32 as=0 ps=0 
M1366 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/an 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/ai gnd nfet w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1367 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/bn 3seg_0/firseg_0/3_bitmux_0/o1 gnd gnd nfet w=6 l=2
+ ad=42 pd=26 as=0 ps=0 
M1368 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/mux_0/a1 vdd vdd pfet w=24 l=2
+ ad=168 pd=64 as=0 ps=0 
M1369 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/a1 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1370 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/mux_0/a1 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1371 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/a1 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1372 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/mux_0/a1 vdd pfet w=27 l=2
+ ad=424 pd=138 as=530 ps=208 
M1373 3seg_0/2seg_0/totdiff3_0/mux_0/a1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn vdd pfet w=27 l=2
+ ad=0 pd=0 as=0 ps=0 
M1374 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/mux_0/a1 vdd pfet w=27 l=2
+ ad=440 pd=142 as=0 ps=0 
M1375 3seg_0/2seg_0/totdiff3_0/mux_0/a1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn vdd pfet w=27 l=2
+ ad=0 pd=0 as=0 ps=0 
M1376 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c vdd vdd pfet w=26 l=2
+ ad=0 pd=0 as=0 ps=0 
M1377 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn vdd pfet w=26 l=2
+ ad=0 pd=0 as=0 ps=0 
M1378 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/iz vdd vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1379 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1380 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/bn vdd pfet w=28 l=2
+ ad=224 pd=72 as=272 ps=122 
M1381 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/iz vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1382 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1383 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/bn 3seg_0/firseg_0/3_bitmux_0/o1 vdd vdd pfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1384 vdd 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/bn vdd pfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1385 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/a_11_12# 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn gnd gnd nfet w=12 l=2
+ ad=60 pd=34 as=0 ps=0 
M1386 3seg_0/2seg_0/totdiff3_0/mux_0/a1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/a_11_12# gnd nfet w=12 l=2
+ ad=208 pd=84 as=0 ps=0 
M1387 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/a_28_12# 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/mux_0/a1 gnd nfet w=12 l=2
+ ad=60 pd=34 as=0 ps=0 
M1388 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/a_28_12# gnd nfet w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1389 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/iz gnd gnd nfet w=14 l=2
+ ad=224 pd=88 as=0 ps=0 
M1390 3seg_0/2seg_0/totdiff3_0/mux_0/a1 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn gnd nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1391 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c 3seg_0/2seg_0/totdiff3_0/mux_0/a1 gnd nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1392 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn gnd nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1393 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c gnd gnd nfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1394 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn gnd nfet w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1395 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/a_115_7# 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1396 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/a_115_7# gnd nfet w=13 l=2
+ ad=104 pd=42 as=0 ps=0 
M1397 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/iz gnd nfet w=13 l=2
+ ad=114 pd=52 as=0 ps=0 
M1398 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a gnd nfet w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1399 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/bn 3seg_0/firseg_0/3_bitmux_0/o1 gnd gnd nfet w=11 l=2
+ ad=67 pd=36 as=0 ps=0 
M1400 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/in_2c vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1401 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1402 vdd vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1403 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/in_2c gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1404 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a_24_13# 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1405 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/zn vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1406 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/mux_0/b0 vdd pfet w=20 l=2
+ ad=320 pd=112 as=398 ps=164 
M1407 3seg_0/2seg_0/totdiff3_0/mux_0/b0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1408 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/mux_0/b0 vdd pfet w=20 l=2
+ ad=320 pd=112 as=0 ps=0 
M1409 3seg_0/2seg_0/totdiff3_0/mux_0/b0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1410 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn vdd vdd vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1411 vdd vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1412 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a vdd vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1413 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1414 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/a_13_13# 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1415 3seg_0/2seg_0/totdiff3_0/mux_0/b0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/a_13_13# gnd nfet w=13 l=2
+ ad=264 pd=98 as=0 ps=0 
M1416 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/a_30_13# 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/mux_0/b0 gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1417 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/a_30_13# gnd nfet w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1418 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn vdd gnd gnd nfet w=10 l=2
+ ad=130 pd=56 as=0 ps=0 
M1419 3seg_0/2seg_0/totdiff3_0/mux_0/b0 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn gnd nfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1420 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an vdd 3seg_0/2seg_0/totdiff3_0/mux_0/b0 gnd nfet w=20 l=2
+ ad=130 pd=56 as=0 ps=0 
M1421 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1422 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1423 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1424 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/a_31_39# 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/z vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1425 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/z 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1426 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/a_48_39# 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/z 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1427 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/z 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1428 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1429 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/z gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1430 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/z 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1431 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1432 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1433 vdd 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1434 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1435 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a_24_13# 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1436 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/zn 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1437 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1438 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/zn gnd vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1439 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/b 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1440 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1441 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/a_24_13# gnd gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1442 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/b 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1443 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/b vdd pfet w=12 l=2
+ ad=0 pd=0 as=72 ps=38 
M1444 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/an 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z vdd vdd pfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1445 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/an vdd pfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1446 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/ai 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/zn vdd pfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1447 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/an 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/ai vdd pfet w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1448 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/bn 3seg_0/firseg_0/3_bitmux_0/o0 vdd vdd pfet w=12 l=2
+ ad=72 pd=38 as=0 ps=0 
M1449 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/b gnd nfet w=6 l=2
+ ad=0 pd=0 as=42 ps=26 
M1450 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/an 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z gnd gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1451 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/zn 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/an gnd nfet w=6 l=2
+ ad=48 pd=28 as=0 ps=0 
M1452 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/ai 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/zn gnd nfet w=6 l=2
+ ad=57 pd=32 as=0 ps=0 
M1453 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/an 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/ai gnd nfet w=6 l=2
+ ad=0 pd=0 as=0 ps=0 
M1454 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/bn 3seg_0/firseg_0/3_bitmux_0/o0 gnd gnd nfet w=6 l=2
+ ad=42 pd=26 as=0 ps=0 
M1455 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/mux_0/a0 vdd vdd pfet w=24 l=2
+ ad=168 pd=64 as=0 ps=0 
M1456 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/a0 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1457 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/mux_0/a0 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1458 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/a0 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1459 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/mux_0/a0 vdd pfet w=27 l=2
+ ad=424 pd=138 as=530 ps=208 
M1460 3seg_0/2seg_0/totdiff3_0/mux_0/a0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn vdd pfet w=27 l=2
+ ad=0 pd=0 as=0 ps=0 
M1461 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/mux_0/a0 vdd pfet w=27 l=2
+ ad=440 pd=142 as=0 ps=0 
M1462 3seg_0/2seg_0/totdiff3_0/mux_0/a0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn vdd pfet w=27 l=2
+ ad=0 pd=0 as=0 ps=0 
M1463 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn gnd vdd vdd pfet w=26 l=2
+ ad=0 pd=0 as=0 ps=0 
M1464 vdd gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn vdd pfet w=26 l=2
+ ad=0 pd=0 as=0 ps=0 
M1465 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/iz vdd vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1466 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1467 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/bn vdd pfet w=28 l=2
+ ad=224 pd=72 as=272 ps=122 
M1468 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/iz vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1469 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1470 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/bn 3seg_0/firseg_0/3_bitmux_0/o0 vdd vdd pfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1471 vdd 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/bn vdd pfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1472 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/a_11_12# 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn gnd gnd nfet w=12 l=2
+ ad=60 pd=34 as=0 ps=0 
M1473 3seg_0/2seg_0/totdiff3_0/mux_0/a0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/a_11_12# gnd nfet w=12 l=2
+ ad=208 pd=84 as=0 ps=0 
M1474 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/a_28_12# 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/mux_0/a0 gnd nfet w=12 l=2
+ ad=60 pd=34 as=0 ps=0 
M1475 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/a_28_12# gnd nfet w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1476 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/iz gnd gnd nfet w=14 l=2
+ ad=224 pd=88 as=0 ps=0 
M1477 3seg_0/2seg_0/totdiff3_0/mux_0/a0 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn gnd nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1478 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn gnd 3seg_0/2seg_0/totdiff3_0/mux_0/a0 gnd nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1479 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn gnd nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1480 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn gnd gnd gnd nfet w=12 l=2
+ ad=96 pd=40 as=0 ps=0 
M1481 gnd gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn gnd nfet w=12 l=2
+ ad=0 pd=0 as=0 ps=0 
M1482 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/a_115_7# 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1483 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/a_115_7# gnd nfet w=13 l=2
+ ad=104 pd=42 as=0 ps=0 
M1484 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/iz gnd nfet w=13 l=2
+ ad=114 pd=52 as=0 ps=0 
M1485 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a gnd nfet w=13 l=2
+ ad=0 pd=0 as=0 ps=0 
M1486 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/bn 3seg_0/firseg_0/3_bitmux_0/o0 gnd gnd nfet w=11 l=2
+ ad=67 pd=36 as=0 ps=0 
M1487 vdd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/zn 3seg_0/firseg_0/3_bitmux_0/o2 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# pfet w=18 l=2
+ ad=0 pd=0 as=102 ps=50 
M1488 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/a_21_50# 3seg_0/firseg_0/decoder_0/b2 vdd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1489 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/zn 3seg_0/firseg_0/out 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/a_21_50# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=128 pd=48 as=0 ps=0 
M1490 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/a_38_50# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/sn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/zn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1491 vdd decoder_0/b2 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/a_38_50# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1492 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/sn 3seg_0/firseg_0/out vdd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# pfet w=8 l=2
+ ad=52 pd=30 as=0 ps=0 
M1493 gnd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/zn 3seg_0/firseg_0/3_bitmux_0/o2 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# nfet w=9 l=2
+ ad=0 pd=0 as=57 ps=32 
M1494 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/a_21_12# 3seg_0/firseg_0/decoder_0/b2 gnd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# nfet w=8 l=2
+ ad=40 pd=26 as=0 ps=0 
M1495 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/zn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/sn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/a_21_12# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# nfet w=8 l=2
+ ad=64 pd=32 as=0 ps=0 
M1496 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/a_38_12# 3seg_0/firseg_0/out 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/zn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# nfet w=8 l=2
+ ad=40 pd=26 as=0 ps=0 
M1497 gnd decoder_0/b2 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/a_38_12# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1498 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/sn 3seg_0/firseg_0/out gnd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# nfet w=6 l=2
+ ad=42 pd=26 as=0 ps=0 
M1499 vdd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/zn 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# pfet w=18 l=2
+ ad=0 pd=0 as=102 ps=50 
M1500 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/a_21_50# 3seg_0/firseg_0/decoder_0/b1 vdd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1501 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/zn 3seg_0/firseg_0/out 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/a_21_50# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=128 pd=48 as=0 ps=0 
M1502 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/a_38_50# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/sn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/zn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1503 vdd decoder_0/b1 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/a_38_50# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1504 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/sn 3seg_0/firseg_0/out vdd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# pfet w=8 l=2
+ ad=52 pd=30 as=0 ps=0 
M1505 gnd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/zn 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# nfet w=9 l=2
+ ad=0 pd=0 as=57 ps=32 
M1506 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/a_21_12# 3seg_0/firseg_0/decoder_0/b1 gnd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=40 pd=26 as=0 ps=0 
M1507 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/zn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/sn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/a_21_12# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=64 pd=32 as=0 ps=0 
M1508 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/a_38_12# 3seg_0/firseg_0/out 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/zn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=40 pd=26 as=0 ps=0 
M1509 gnd decoder_0/b1 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/a_38_12# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1510 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/sn 3seg_0/firseg_0/out gnd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# nfet w=6 l=2
+ ad=42 pd=26 as=0 ps=0 
M1511 vdd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/zn 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# pfet w=18 l=2
+ ad=0 pd=0 as=102 ps=50 
M1512 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/a_21_50# 3seg_0/firseg_0/decoder_0/b0 vdd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1513 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/zn 3seg_0/firseg_0/out 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/a_21_50# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# pfet w=16 l=2
+ ad=128 pd=48 as=0 ps=0 
M1514 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/a_38_50# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/sn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/zn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1515 vdd decoder_0/b0 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/a_38_50# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1516 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/sn 3seg_0/firseg_0/out vdd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# pfet w=8 l=2
+ ad=52 pd=30 as=0 ps=0 
M1517 gnd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/zn 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# nfet w=9 l=2
+ ad=0 pd=0 as=57 ps=32 
M1518 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/a_21_12# 3seg_0/firseg_0/decoder_0/b0 gnd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=40 pd=26 as=0 ps=0 
M1519 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/zn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/sn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/a_21_12# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=64 pd=32 as=0 ps=0 
M1520 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/a_38_12# 3seg_0/firseg_0/out 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/zn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=40 pd=26 as=0 ps=0 
M1521 gnd decoder_0/b0 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/a_38_12# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1522 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/sn 3seg_0/firseg_0/out gnd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# nfet w=6 l=2
+ ad=42 pd=26 as=0 ps=0 
M1523 3seg_0/firseg_0/out 3seg_0/firseg_0/comp_0/nr3v0x2_0/z vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=14 l=2
+ ad=392 pd=120 as=0 ps=0 
M1524 vdd 3seg_0/firseg_0/comp_0/nr3v0x2_0/z 3seg_0/firseg_0/out 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1525 3seg_0/firseg_0/out 3seg_0/firseg_0/comp_0/nd3v0x2_0/c vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1526 vdd 3seg_0/firseg_0/comp_0/nd3v0x2_0/a 3seg_0/firseg_0/out 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1527 3seg_0/firseg_0/comp_0/nd3v0x2_0/a_14_12# 3seg_0/firseg_0/comp_0/nd3v0x2_0/a gnd gnd nfet w=14 l=2
+ ad=70 pd=38 as=0 ps=0 
M1528 3seg_0/firseg_0/comp_0/nd3v0x2_0/a_21_12# 3seg_0/firseg_0/comp_0/nr3v0x2_0/z 3seg_0/firseg_0/comp_0/nd3v0x2_0/a_14_12# gnd nfet w=14 l=2
+ ad=70 pd=38 as=0 ps=0 
M1529 3seg_0/firseg_0/out 3seg_0/firseg_0/comp_0/nd3v0x2_0/c 3seg_0/firseg_0/comp_0/nd3v0x2_0/a_21_12# gnd nfet w=14 l=2
+ ad=112 pd=44 as=0 ps=0 
M1530 3seg_0/firseg_0/comp_0/nd3v0x2_0/a_38_12# 3seg_0/firseg_0/comp_0/nd3v0x2_0/c 3seg_0/firseg_0/out gnd nfet w=14 l=2
+ ad=70 pd=38 as=0 ps=0 
M1531 3seg_0/firseg_0/comp_0/nd3v0x2_0/a_45_12# 3seg_0/firseg_0/comp_0/nr3v0x2_0/z 3seg_0/firseg_0/comp_0/nd3v0x2_0/a_38_12# gnd nfet w=14 l=2
+ ad=70 pd=38 as=0 ps=0 
M1532 gnd 3seg_0/firseg_0/comp_0/nd3v0x2_0/a 3seg_0/firseg_0/comp_0/nd3v0x2_0/a_45_12# gnd nfet w=14 l=2
+ ad=0 pd=0 as=0 ps=0 
M1533 vdd 3seg_0/firseg_0/comp_0/an3v0x2_1/zn 3seg_0/firseg_0/comp_0/nr2v0x2_1/a 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1534 3seg_0/firseg_0/comp_0/an3v0x2_1/zn 3seg_0/firseg_0/comp_0/an3v0x2_1/a vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=17 l=2
+ ad=233 pd=98 as=0 ps=0 
M1535 vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/b 3seg_0/firseg_0/comp_0/an3v0x2_1/zn 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=17 l=2
+ ad=0 pd=0 as=0 ps=0 
M1536 3seg_0/firseg_0/comp_0/an3v0x2_1/zn 3seg_0/firseg_0/decoder_0/b2 vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=17 l=2
+ ad=0 pd=0 as=0 ps=0 
M1537 gnd 3seg_0/firseg_0/comp_0/an3v0x2_1/zn 3seg_0/firseg_0/comp_0/nr2v0x2_1/a gnd nfet w=14 l=2
+ ad=0 pd=0 as=82 ps=42 
M1538 3seg_0/firseg_0/comp_0/an3v0x2_1/a_24_8# 3seg_0/firseg_0/comp_0/an3v0x2_1/a gnd gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1539 3seg_0/firseg_0/comp_0/an3v0x2_1/a_31_8# 3seg_0/firseg_0/comp_0/an3v0x2_2/b 3seg_0/firseg_0/comp_0/an3v0x2_1/a_24_8# gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1540 3seg_0/firseg_0/comp_0/an3v0x2_1/zn 3seg_0/firseg_0/decoder_0/b2 3seg_0/firseg_0/comp_0/an3v0x2_1/a_31_8# gnd nfet w=17 l=2
+ ad=97 pd=48 as=0 ps=0 
M1541 3seg_0/firseg_0/comp_0/nr3v0x2_0/a_13_39# 3seg_0/firseg_0/comp_0/an3v0x2_2/z 3seg_0/firseg_0/comp_0/nr3v0x2_0/z 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=27 l=2
+ ad=135 pd=64 as=377 ps=138 
M1542 3seg_0/firseg_0/comp_0/nr3v0x2_0/a_20_39# 3seg_0/firseg_0/comp_0/an3v0x2_0/z 3seg_0/firseg_0/comp_0/nr3v0x2_0/a_13_39# 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=27 l=2
+ ad=135 pd=64 as=0 ps=0 
M1543 vdd 3seg_0/firseg_0/comp_0/nr3v0x2_0/a 3seg_0/firseg_0/comp_0/nr3v0x2_0/a_20_39# 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=27 l=2
+ ad=0 pd=0 as=0 ps=0 
M1544 3seg_0/firseg_0/comp_0/nr3v0x2_0/a_37_39# 3seg_0/firseg_0/comp_0/nr3v0x2_0/a vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=27 l=2
+ ad=135 pd=64 as=0 ps=0 
M1545 3seg_0/firseg_0/comp_0/nr3v0x2_0/a_44_39# 3seg_0/firseg_0/comp_0/an3v0x2_0/z 3seg_0/firseg_0/comp_0/nr3v0x2_0/a_37_39# 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=27 l=2
+ ad=135 pd=64 as=0 ps=0 
M1546 3seg_0/firseg_0/comp_0/nr3v0x2_0/z 3seg_0/firseg_0/comp_0/an3v0x2_2/z 3seg_0/firseg_0/comp_0/nr3v0x2_0/a_44_39# 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=27 l=2
+ ad=0 pd=0 as=0 ps=0 
M1547 3seg_0/firseg_0/comp_0/nr3v0x2_0/a_61_39# 3seg_0/firseg_0/comp_0/an3v0x2_2/z 3seg_0/firseg_0/comp_0/nr3v0x2_0/z 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=27 l=2
+ ad=135 pd=64 as=0 ps=0 
M1548 3seg_0/firseg_0/comp_0/nr3v0x2_0/a_68_39# 3seg_0/firseg_0/comp_0/an3v0x2_0/z 3seg_0/firseg_0/comp_0/nr3v0x2_0/a_61_39# 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=27 l=2
+ ad=135 pd=64 as=0 ps=0 
M1549 vdd 3seg_0/firseg_0/comp_0/nr3v0x2_0/a 3seg_0/firseg_0/comp_0/nr3v0x2_0/a_68_39# 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=27 l=2
+ ad=0 pd=0 as=0 ps=0 
M1550 gnd 3seg_0/firseg_0/comp_0/an3v0x2_2/z 3seg_0/firseg_0/comp_0/nr3v0x2_0/z gnd nfet w=15 l=2
+ ad=0 pd=0 as=207 ps=90 
M1551 3seg_0/firseg_0/comp_0/nr3v0x2_0/z 3seg_0/firseg_0/comp_0/an3v0x2_0/z gnd gnd nfet w=15 l=2
+ ad=0 pd=0 as=0 ps=0 
M1552 gnd 3seg_0/firseg_0/comp_0/nr3v0x2_0/a 3seg_0/firseg_0/comp_0/nr3v0x2_0/z gnd nfet w=15 l=2
+ ad=0 pd=0 as=0 ps=0 
M1553 vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/zn 3seg_0/firseg_0/comp_0/an3v0x2_2/z 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1554 3seg_0/firseg_0/comp_0/an3v0x2_2/zn 3seg_0/firseg_0/decoder_0/b0 vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=17 l=2
+ ad=233 pd=98 as=0 ps=0 
M1555 vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/b 3seg_0/firseg_0/comp_0/an3v0x2_2/zn 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=17 l=2
+ ad=0 pd=0 as=0 ps=0 
M1556 3seg_0/firseg_0/comp_0/an3v0x2_2/zn 3seg_0/firseg_0/decoder_0/b2 vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# pfet w=17 l=2
+ ad=0 pd=0 as=0 ps=0 
M1557 gnd 3seg_0/firseg_0/comp_0/an3v0x2_2/zn 3seg_0/firseg_0/comp_0/an3v0x2_2/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=82 ps=42 
M1558 3seg_0/firseg_0/comp_0/an3v0x2_2/a_24_8# 3seg_0/firseg_0/decoder_0/b0 gnd gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1559 3seg_0/firseg_0/comp_0/an3v0x2_2/a_31_8# 3seg_0/firseg_0/comp_0/an3v0x2_2/b 3seg_0/firseg_0/comp_0/an3v0x2_2/a_24_8# gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1560 3seg_0/firseg_0/comp_0/an3v0x2_2/zn 3seg_0/firseg_0/decoder_0/b2 3seg_0/firseg_0/comp_0/an3v0x2_2/a_31_8# gnd nfet w=17 l=2
+ ad=97 pd=48 as=0 ps=0 
M1561 3seg_0/firseg_0/comp_0/nr2v0x2_1/a_11_39# 3seg_0/firseg_0/comp_0/nr2v0x2_1/a vdd vdd pfet w=27 l=2
+ ad=135 pd=64 as=0 ps=0 
M1562 3seg_0/firseg_0/comp_0/nd3v0x2_0/c 3seg_0/firseg_0/comp_0/an3v0x2_3/z 3seg_0/firseg_0/comp_0/nr2v0x2_1/a_11_39# vdd pfet w=27 l=2
+ ad=216 pd=70 as=0 ps=0 
M1563 3seg_0/firseg_0/comp_0/nr2v0x2_1/a_28_39# 3seg_0/firseg_0/comp_0/an3v0x2_3/z 3seg_0/firseg_0/comp_0/nd3v0x2_0/c vdd pfet w=27 l=2
+ ad=135 pd=64 as=0 ps=0 
M1564 vdd 3seg_0/firseg_0/comp_0/nr2v0x2_1/a 3seg_0/firseg_0/comp_0/nr2v0x2_1/a_28_39# vdd pfet w=27 l=2
+ ad=0 pd=0 as=0 ps=0 
M1565 3seg_0/firseg_0/comp_0/nd3v0x2_0/c 3seg_0/firseg_0/comp_0/nr2v0x2_1/a gnd gnd nfet w=15 l=2
+ ad=120 pd=46 as=0 ps=0 
M1566 gnd 3seg_0/firseg_0/comp_0/an3v0x2_3/z 3seg_0/firseg_0/comp_0/nd3v0x2_0/c gnd nfet w=15 l=2
+ ad=0 pd=0 as=0 ps=0 
M1567 vdd 3seg_0/firseg_0/comp_0/an3v0x2_3/zn 3seg_0/firseg_0/comp_0/an3v0x2_3/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1568 3seg_0/firseg_0/comp_0/an3v0x2_3/zn 3seg_0/firseg_0/comp_0/an2v0x2_0/b vdd vdd pfet w=17 l=2
+ ad=233 pd=98 as=0 ps=0 
M1569 vdd 3seg_0/firseg_0/decoder_0/b1 3seg_0/firseg_0/comp_0/an3v0x2_3/zn vdd pfet w=17 l=2
+ ad=0 pd=0 as=0 ps=0 
M1570 3seg_0/firseg_0/comp_0/an3v0x2_3/zn 3seg_0/firseg_0/decoder_0/b0 vdd vdd pfet w=17 l=2
+ ad=0 pd=0 as=0 ps=0 
M1571 gnd 3seg_0/firseg_0/comp_0/an3v0x2_3/zn 3seg_0/firseg_0/comp_0/an3v0x2_3/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=82 ps=42 
M1572 3seg_0/firseg_0/comp_0/an3v0x2_3/a_24_8# 3seg_0/firseg_0/comp_0/an2v0x2_0/b gnd gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1573 3seg_0/firseg_0/comp_0/an3v0x2_3/a_31_8# 3seg_0/firseg_0/decoder_0/b1 3seg_0/firseg_0/comp_0/an3v0x2_3/a_24_8# gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1574 3seg_0/firseg_0/comp_0/an3v0x2_3/zn 3seg_0/firseg_0/decoder_0/b0 3seg_0/firseg_0/comp_0/an3v0x2_3/a_31_8# gnd nfet w=17 l=2
+ ad=97 pd=48 as=0 ps=0 
M1575 vdd 3seg_0/firseg_0/comp_0/an3v0x2_0/zn 3seg_0/firseg_0/comp_0/an3v0x2_0/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1576 3seg_0/firseg_0/comp_0/an3v0x2_0/zn 3seg_0/firseg_0/comp_0/an3v0x2_1/a vdd vdd pfet w=17 l=2
+ ad=233 pd=98 as=0 ps=0 
M1577 vdd 3seg_0/firseg_0/decoder_0/b1 3seg_0/firseg_0/comp_0/an3v0x2_0/zn vdd pfet w=17 l=2
+ ad=0 pd=0 as=0 ps=0 
M1578 3seg_0/firseg_0/comp_0/an3v0x2_0/zn 3seg_0/firseg_0/comp_0/an2v0x2_0/b vdd vdd pfet w=17 l=2
+ ad=0 pd=0 as=0 ps=0 
M1579 gnd 3seg_0/firseg_0/comp_0/an3v0x2_0/zn 3seg_0/firseg_0/comp_0/an3v0x2_0/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=82 ps=42 
M1580 3seg_0/firseg_0/comp_0/an3v0x2_0/a_24_8# 3seg_0/firseg_0/comp_0/an3v0x2_1/a gnd gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1581 3seg_0/firseg_0/comp_0/an3v0x2_0/a_31_8# 3seg_0/firseg_0/decoder_0/b1 3seg_0/firseg_0/comp_0/an3v0x2_0/a_24_8# gnd nfet w=17 l=2
+ ad=85 pd=44 as=0 ps=0 
M1582 3seg_0/firseg_0/comp_0/an3v0x2_0/zn 3seg_0/firseg_0/comp_0/an2v0x2_0/b 3seg_0/firseg_0/comp_0/an3v0x2_0/a_31_8# gnd nfet w=17 l=2
+ ad=97 pd=48 as=0 ps=0 
M1583 vdd 3seg_0/firseg_0/comp_0/an2v0x2_0/zn 3seg_0/firseg_0/comp_0/nr3v0x2_0/a vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1584 3seg_0/firseg_0/comp_0/an2v0x2_0/zn 3seg_0/firseg_0/decoder_0/b2 vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1585 vdd 3seg_0/firseg_0/comp_0/an2v0x2_0/b 3seg_0/firseg_0/comp_0/an2v0x2_0/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1586 gnd 3seg_0/firseg_0/comp_0/an2v0x2_0/zn 3seg_0/firseg_0/comp_0/nr3v0x2_0/a gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1587 3seg_0/firseg_0/comp_0/an2v0x2_0/a_24_13# 3seg_0/firseg_0/decoder_0/b2 gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1588 3seg_0/firseg_0/comp_0/an2v0x2_0/zn 3seg_0/firseg_0/comp_0/an2v0x2_0/b 3seg_0/firseg_0/comp_0/an2v0x2_0/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1589 3seg_0/firseg_0/comp_0/nr2v0x2_0/a_11_39# 3seg_0/firseg_0/comp_0/an2v0x2_3/z vdd vdd pfet w=27 l=2
+ ad=135 pd=64 as=0 ps=0 
M1590 3seg_0/firseg_0/comp_0/nd3v0x2_0/a 3seg_0/firseg_0/comp_0/an2v0x2_1/z 3seg_0/firseg_0/comp_0/nr2v0x2_0/a_11_39# vdd pfet w=27 l=2
+ ad=216 pd=70 as=0 ps=0 
M1591 3seg_0/firseg_0/comp_0/nr2v0x2_0/a_28_39# 3seg_0/firseg_0/comp_0/an2v0x2_1/z 3seg_0/firseg_0/comp_0/nd3v0x2_0/a vdd pfet w=27 l=2
+ ad=135 pd=64 as=0 ps=0 
M1592 vdd 3seg_0/firseg_0/comp_0/an2v0x2_3/z 3seg_0/firseg_0/comp_0/nr2v0x2_0/a_28_39# vdd pfet w=27 l=2
+ ad=0 pd=0 as=0 ps=0 
M1593 3seg_0/firseg_0/comp_0/nd3v0x2_0/a 3seg_0/firseg_0/comp_0/an2v0x2_3/z gnd gnd nfet w=15 l=2
+ ad=120 pd=46 as=0 ps=0 
M1594 gnd 3seg_0/firseg_0/comp_0/an2v0x2_1/z 3seg_0/firseg_0/comp_0/nd3v0x2_0/a gnd nfet w=15 l=2
+ ad=0 pd=0 as=0 ps=0 
M1595 vdd 3seg_0/firseg_0/comp_0/or3v0x2_1/zn 3seg_0/firseg_0/comp_0/an2v0x2_3/b vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1596 3seg_0/firseg_0/comp_0/or3v0x2_1/a_24_38# 3seg_0/firseg_0/comp_0/an3v0x2_2/b vdd vdd pfet w=22 l=2
+ ad=110 pd=54 as=0 ps=0 
M1597 3seg_0/firseg_0/comp_0/or3v0x2_1/a_31_38# 3seg_0/firseg_0/comp_0/an3v0x2_1/a 3seg_0/firseg_0/comp_0/or3v0x2_1/a_24_38# vdd pfet w=22 l=2
+ ad=110 pd=54 as=0 ps=0 
M1598 3seg_0/firseg_0/comp_0/or3v0x2_1/zn 3seg_0/firseg_0/decoder_0/b0 3seg_0/firseg_0/comp_0/or3v0x2_1/a_31_38# vdd pfet w=22 l=2
+ ad=167 pd=60 as=0 ps=0 
M1599 3seg_0/firseg_0/comp_0/or3v0x2_1/a_48_38# 3seg_0/firseg_0/decoder_0/b0 3seg_0/firseg_0/comp_0/or3v0x2_1/zn vdd pfet w=19 l=2
+ ad=95 pd=48 as=0 ps=0 
M1600 3seg_0/firseg_0/comp_0/or3v0x2_1/a_55_38# 3seg_0/firseg_0/comp_0/an3v0x2_1/a 3seg_0/firseg_0/comp_0/or3v0x2_1/a_48_38# vdd pfet w=19 l=2
+ ad=95 pd=48 as=0 ps=0 
M1601 vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/b 3seg_0/firseg_0/comp_0/or3v0x2_1/a_55_38# vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1602 gnd 3seg_0/firseg_0/comp_0/or3v0x2_1/zn 3seg_0/firseg_0/comp_0/an2v0x2_3/b gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1603 3seg_0/firseg_0/comp_0/or3v0x2_1/zn 3seg_0/firseg_0/comp_0/an3v0x2_2/b gnd gnd nfet w=8 l=2
+ ad=116 pd=62 as=0 ps=0 
M1604 gnd 3seg_0/firseg_0/comp_0/an3v0x2_1/a 3seg_0/firseg_0/comp_0/or3v0x2_1/zn gnd nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1605 3seg_0/firseg_0/comp_0/or3v0x2_1/zn 3seg_0/firseg_0/decoder_0/b0 gnd gnd nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1606 vdd 3seg_0/firseg_0/comp_0/an2v0x2_1/zn 3seg_0/firseg_0/comp_0/an2v0x2_1/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1607 3seg_0/firseg_0/comp_0/an2v0x2_1/zn 3seg_0/firseg_0/comp_0/an2v0x2_4/z vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1608 vdd 3seg_0/firseg_0/comp_0/an2v0x2_1/b 3seg_0/firseg_0/comp_0/an2v0x2_1/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1609 gnd 3seg_0/firseg_0/comp_0/an2v0x2_1/zn 3seg_0/firseg_0/comp_0/an2v0x2_1/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1610 3seg_0/firseg_0/comp_0/an2v0x2_1/a_24_13# 3seg_0/firseg_0/comp_0/an2v0x2_4/z gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1611 3seg_0/firseg_0/comp_0/an2v0x2_1/zn 3seg_0/firseg_0/comp_0/an2v0x2_1/b 3seg_0/firseg_0/comp_0/an2v0x2_1/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1612 vdd 3seg_0/firseg_0/comp_0/an2v0x2_4/zn 3seg_0/firseg_0/comp_0/an2v0x2_4/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1613 3seg_0/firseg_0/comp_0/an2v0x2_4/zn 3seg_0/firseg_0/comp_0/an2v0x2_0/b vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1614 vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/b 3seg_0/firseg_0/comp_0/an2v0x2_4/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1615 gnd 3seg_0/firseg_0/comp_0/an2v0x2_4/zn 3seg_0/firseg_0/comp_0/an2v0x2_4/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1616 3seg_0/firseg_0/comp_0/an2v0x2_4/a_24_13# 3seg_0/firseg_0/comp_0/an2v0x2_0/b gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1617 3seg_0/firseg_0/comp_0/an2v0x2_4/zn 3seg_0/firseg_0/comp_0/an3v0x2_2/b 3seg_0/firseg_0/comp_0/an2v0x2_4/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1618 3seg_0/firseg_0/comp_0/an3v0x2_2/b decoder_0/b1 vdd vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1619 vdd decoder_0/b1 3seg_0/firseg_0/comp_0/an3v0x2_2/b vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1620 3seg_0/firseg_0/comp_0/an3v0x2_2/b decoder_0/b1 gnd gnd nfet w=17 l=2
+ ad=118 pd=50 as=0 ps=0 
M1621 gnd decoder_0/b1 3seg_0/firseg_0/comp_0/an3v0x2_2/b gnd nfet w=11 l=2
+ ad=0 pd=0 as=0 ps=0 
M1622 vdd 3seg_0/firseg_0/comp_0/an2v0x2_3/zn 3seg_0/firseg_0/comp_0/an2v0x2_3/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1623 3seg_0/firseg_0/comp_0/an2v0x2_3/zn 3seg_0/firseg_0/comp_0/an2v0x2_2/z vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1624 vdd 3seg_0/firseg_0/comp_0/an2v0x2_3/b 3seg_0/firseg_0/comp_0/an2v0x2_3/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1625 gnd 3seg_0/firseg_0/comp_0/an2v0x2_3/zn 3seg_0/firseg_0/comp_0/an2v0x2_3/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1626 3seg_0/firseg_0/comp_0/an2v0x2_3/a_24_13# 3seg_0/firseg_0/comp_0/an2v0x2_2/z gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1627 3seg_0/firseg_0/comp_0/an2v0x2_3/zn 3seg_0/firseg_0/comp_0/an2v0x2_3/b 3seg_0/firseg_0/comp_0/an2v0x2_3/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1628 vdd 3seg_0/firseg_0/comp_0/an2v0x2_2/zn 3seg_0/firseg_0/comp_0/an2v0x2_2/z vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1629 3seg_0/firseg_0/comp_0/an2v0x2_2/zn 3seg_0/firseg_0/decoder_0/b2 vdd vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1630 vdd 3seg_0/firseg_0/decoder_0/b1 3seg_0/firseg_0/comp_0/an2v0x2_2/zn vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1631 gnd 3seg_0/firseg_0/comp_0/an2v0x2_2/zn 3seg_0/firseg_0/comp_0/an2v0x2_2/z gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1632 3seg_0/firseg_0/comp_0/an2v0x2_2/a_24_13# 3seg_0/firseg_0/decoder_0/b2 gnd gnd nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1633 3seg_0/firseg_0/comp_0/an2v0x2_2/zn 3seg_0/firseg_0/decoder_0/b1 3seg_0/firseg_0/comp_0/an2v0x2_2/a_24_13# gnd nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1634 vdd 3seg_0/firseg_0/comp_0/or3v0x2_0/zn 3seg_0/firseg_0/comp_0/an2v0x2_1/b vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1635 3seg_0/firseg_0/comp_0/or3v0x2_0/a_24_38# 3seg_0/firseg_0/decoder_0/b1 vdd vdd pfet w=22 l=2
+ ad=110 pd=54 as=0 ps=0 
M1636 3seg_0/firseg_0/comp_0/or3v0x2_0/a_31_38# 3seg_0/firseg_0/decoder_0/b0 3seg_0/firseg_0/comp_0/or3v0x2_0/a_24_38# vdd pfet w=22 l=2
+ ad=110 pd=54 as=0 ps=0 
M1637 3seg_0/firseg_0/comp_0/or3v0x2_0/zn 3seg_0/firseg_0/comp_0/an3v0x2_1/a 3seg_0/firseg_0/comp_0/or3v0x2_0/a_31_38# vdd pfet w=22 l=2
+ ad=167 pd=60 as=0 ps=0 
M1638 3seg_0/firseg_0/comp_0/or3v0x2_0/a_48_38# 3seg_0/firseg_0/comp_0/an3v0x2_1/a 3seg_0/firseg_0/comp_0/or3v0x2_0/zn vdd pfet w=19 l=2
+ ad=95 pd=48 as=0 ps=0 
M1639 3seg_0/firseg_0/comp_0/or3v0x2_0/a_55_38# 3seg_0/firseg_0/decoder_0/b0 3seg_0/firseg_0/comp_0/or3v0x2_0/a_48_38# vdd pfet w=19 l=2
+ ad=95 pd=48 as=0 ps=0 
M1640 vdd 3seg_0/firseg_0/decoder_0/b1 3seg_0/firseg_0/comp_0/or3v0x2_0/a_55_38# vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1641 gnd 3seg_0/firseg_0/comp_0/or3v0x2_0/zn 3seg_0/firseg_0/comp_0/an2v0x2_1/b gnd nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1642 3seg_0/firseg_0/comp_0/or3v0x2_0/zn 3seg_0/firseg_0/decoder_0/b1 gnd gnd nfet w=8 l=2
+ ad=116 pd=62 as=0 ps=0 
M1643 gnd 3seg_0/firseg_0/decoder_0/b0 3seg_0/firseg_0/comp_0/or3v0x2_0/zn gnd nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1644 3seg_0/firseg_0/comp_0/or3v0x2_0/zn 3seg_0/firseg_0/comp_0/an3v0x2_1/a gnd gnd nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1645 3seg_0/firseg_0/comp_0/an3v0x2_1/a decoder_0/b0 vdd vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1646 vdd decoder_0/b0 3seg_0/firseg_0/comp_0/an3v0x2_1/a vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1647 3seg_0/firseg_0/comp_0/an3v0x2_1/a decoder_0/b0 gnd gnd nfet w=17 l=2
+ ad=118 pd=50 as=0 ps=0 
M1648 gnd decoder_0/b0 3seg_0/firseg_0/comp_0/an3v0x2_1/a gnd nfet w=11 l=2
+ ad=0 pd=0 as=0 ps=0 
M1649 3seg_0/firseg_0/comp_0/an2v0x2_0/b decoder_0/b2 vdd vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1650 vdd decoder_0/b2 3seg_0/firseg_0/comp_0/an2v0x2_0/b vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1651 3seg_0/firseg_0/comp_0/an2v0x2_0/b decoder_0/b2 gnd gnd nfet w=17 l=2
+ ad=118 pd=50 as=0 ps=0 
M1652 gnd decoder_0/b2 3seg_0/firseg_0/comp_0/an2v0x2_0/b gnd nfet w=11 l=2
+ ad=0 pd=0 as=0 ps=0 
M1653 3seg_0/firseg_0/decoder_0/b2 3seg_0/firseg_0/decoder_0/or2v0x3_8/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1654 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_8/zn 3seg_0/firseg_0/decoder_0/b2 vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1655 3seg_0/firseg_0/decoder_0/or2v0x3_8/a_31_39# 3seg_0/firseg_0/decoder_0/d6 vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1656 3seg_0/firseg_0/decoder_0/or2v0x3_8/zn 3seg_0/firseg_0/decoder_0/or2v0x3_7/z 3seg_0/firseg_0/decoder_0/or2v0x3_8/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1657 3seg_0/firseg_0/decoder_0/or2v0x3_8/a_48_39# 3seg_0/firseg_0/decoder_0/or2v0x3_7/z 3seg_0/firseg_0/decoder_0/or2v0x3_8/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1658 vdd 3seg_0/firseg_0/decoder_0/d6 3seg_0/firseg_0/decoder_0/or2v0x3_8/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1659 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_8/zn 3seg_0/firseg_0/decoder_0/b2 gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1660 3seg_0/firseg_0/decoder_0/or2v0x3_8/zn 3seg_0/firseg_0/decoder_0/d6 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1661 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_7/z 3seg_0/firseg_0/decoder_0/or2v0x3_8/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1662 3seg_0/firseg_0/decoder_0/or2v0x3_7/z 3seg_0/firseg_0/decoder_0/or2v0x3_7/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1663 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_7/zn 3seg_0/firseg_0/decoder_0/or2v0x3_7/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1664 3seg_0/firseg_0/decoder_0/or2v0x3_7/a_31_39# 3seg_0/firseg_0/decoder_0/or2v0x3_6/z vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1665 3seg_0/firseg_0/decoder_0/or2v0x3_7/zn 3seg_0/firseg_0/decoder_0/d4 3seg_0/firseg_0/decoder_0/or2v0x3_7/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1666 3seg_0/firseg_0/decoder_0/or2v0x3_7/a_48_39# 3seg_0/firseg_0/decoder_0/d4 3seg_0/firseg_0/decoder_0/or2v0x3_7/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1667 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_6/z 3seg_0/firseg_0/decoder_0/or2v0x3_7/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1668 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_7/zn 3seg_0/firseg_0/decoder_0/or2v0x3_7/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1669 3seg_0/firseg_0/decoder_0/or2v0x3_7/zn 3seg_0/firseg_0/decoder_0/or2v0x3_6/z gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1670 gnd 3seg_0/firseg_0/decoder_0/d4 3seg_0/firseg_0/decoder_0/or2v0x3_7/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1671 3seg_0/firseg_0/decoder_0/or2v0x3_6/z 3seg_0/firseg_0/decoder_0/or2v0x3_6/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1672 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_6/zn 3seg_0/firseg_0/decoder_0/or2v0x3_6/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1673 3seg_0/firseg_0/decoder_0/or2v0x3_6/a_31_39# 3seg_0/firseg_0/decoder_0/d3 vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1674 3seg_0/firseg_0/decoder_0/or2v0x3_6/zn 3seg_0/firseg_0/decoder_0/d5 3seg_0/firseg_0/decoder_0/or2v0x3_6/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1675 3seg_0/firseg_0/decoder_0/or2v0x3_6/a_48_39# 3seg_0/firseg_0/decoder_0/d5 3seg_0/firseg_0/decoder_0/or2v0x3_6/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1676 vdd 3seg_0/firseg_0/decoder_0/d3 3seg_0/firseg_0/decoder_0/or2v0x3_6/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1677 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_6/zn 3seg_0/firseg_0/decoder_0/or2v0x3_6/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1678 3seg_0/firseg_0/decoder_0/or2v0x3_6/zn 3seg_0/firseg_0/decoder_0/d3 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1679 gnd 3seg_0/firseg_0/decoder_0/d5 3seg_0/firseg_0/decoder_0/or2v0x3_6/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1680 3seg_0/firseg_0/decoder_0/b1 3seg_0/firseg_0/decoder_0/or2v0x3_5/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1681 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_5/zn 3seg_0/firseg_0/decoder_0/b1 vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1682 3seg_0/firseg_0/decoder_0/or2v0x3_5/a_31_39# 3seg_0/firseg_0/decoder_0/or2v0x3_4/z vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1683 3seg_0/firseg_0/decoder_0/or2v0x3_5/zn 3seg_0/firseg_0/decoder_0/d6 3seg_0/firseg_0/decoder_0/or2v0x3_5/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1684 3seg_0/firseg_0/decoder_0/or2v0x3_5/a_48_39# 3seg_0/firseg_0/decoder_0/d6 3seg_0/firseg_0/decoder_0/or2v0x3_5/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1685 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_4/z 3seg_0/firseg_0/decoder_0/or2v0x3_5/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1686 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_5/zn 3seg_0/firseg_0/decoder_0/b1 gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1687 3seg_0/firseg_0/decoder_0/or2v0x3_5/zn 3seg_0/firseg_0/decoder_0/or2v0x3_4/z gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1688 gnd 3seg_0/firseg_0/decoder_0/d6 3seg_0/firseg_0/decoder_0/or2v0x3_5/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1689 3seg_0/firseg_0/decoder_0/or2v0x3_4/z 3seg_0/firseg_0/decoder_0/or2v0x3_4/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1690 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_4/zn 3seg_0/firseg_0/decoder_0/or2v0x3_4/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1691 3seg_0/firseg_0/decoder_0/or2v0x3_4/a_31_39# 3seg_0/firseg_0/decoder_0/d1 vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1692 3seg_0/firseg_0/decoder_0/or2v0x3_4/zn 3seg_0/firseg_0/decoder_0/or2v0x3_3/z 3seg_0/firseg_0/decoder_0/or2v0x3_4/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1693 3seg_0/firseg_0/decoder_0/or2v0x3_4/a_48_39# 3seg_0/firseg_0/decoder_0/or2v0x3_3/z 3seg_0/firseg_0/decoder_0/or2v0x3_4/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1694 vdd 3seg_0/firseg_0/decoder_0/d1 3seg_0/firseg_0/decoder_0/or2v0x3_4/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1695 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_4/zn 3seg_0/firseg_0/decoder_0/or2v0x3_4/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1696 3seg_0/firseg_0/decoder_0/or2v0x3_4/zn 3seg_0/firseg_0/decoder_0/d1 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1697 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_3/z 3seg_0/firseg_0/decoder_0/or2v0x3_4/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1698 3seg_0/firseg_0/decoder_0/or2v0x3_3/z 3seg_0/firseg_0/decoder_0/or2v0x3_3/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1699 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_3/zn 3seg_0/firseg_0/decoder_0/or2v0x3_3/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1700 3seg_0/firseg_0/decoder_0/or2v0x3_3/a_31_39# 3seg_0/firseg_0/decoder_0/d5 vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1701 3seg_0/firseg_0/decoder_0/or2v0x3_3/zn 3seg_0/firseg_0/decoder_0/d2 3seg_0/firseg_0/decoder_0/or2v0x3_3/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1702 3seg_0/firseg_0/decoder_0/or2v0x3_3/a_48_39# 3seg_0/firseg_0/decoder_0/d2 3seg_0/firseg_0/decoder_0/or2v0x3_3/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1703 vdd 3seg_0/firseg_0/decoder_0/d5 3seg_0/firseg_0/decoder_0/or2v0x3_3/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1704 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_3/zn 3seg_0/firseg_0/decoder_0/or2v0x3_3/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1705 3seg_0/firseg_0/decoder_0/or2v0x3_3/zn 3seg_0/firseg_0/decoder_0/d5 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1706 gnd 3seg_0/firseg_0/decoder_0/d2 3seg_0/firseg_0/decoder_0/or2v0x3_3/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1707 3seg_0/firseg_0/decoder_0/b0 3seg_0/firseg_0/decoder_0/or2v0x3_2/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1708 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_2/zn 3seg_0/firseg_0/decoder_0/b0 vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1709 3seg_0/firseg_0/decoder_0/or2v0x3_2/a_31_39# 3seg_0/firseg_0/decoder_0/or2v0x3_1/z vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1710 3seg_0/firseg_0/decoder_0/or2v0x3_2/zn 3seg_0/firseg_0/decoder_0/d6 3seg_0/firseg_0/decoder_0/or2v0x3_2/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1711 3seg_0/firseg_0/decoder_0/or2v0x3_2/a_48_39# 3seg_0/firseg_0/decoder_0/d6 3seg_0/firseg_0/decoder_0/or2v0x3_2/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1712 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_1/z 3seg_0/firseg_0/decoder_0/or2v0x3_2/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1713 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_2/zn 3seg_0/firseg_0/decoder_0/b0 gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1714 3seg_0/firseg_0/decoder_0/or2v0x3_2/zn 3seg_0/firseg_0/decoder_0/or2v0x3_1/z gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1715 gnd 3seg_0/firseg_0/decoder_0/d6 3seg_0/firseg_0/decoder_0/or2v0x3_2/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1716 3seg_0/firseg_0/decoder_0/or2v0x3_1/z 3seg_0/firseg_0/decoder_0/or2v0x3_1/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1717 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_1/zn 3seg_0/firseg_0/decoder_0/or2v0x3_1/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1718 3seg_0/firseg_0/decoder_0/or2v0x3_1/a_31_39# 3seg_0/firseg_0/decoder_0/or2v0x3_0/z vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1719 3seg_0/firseg_0/decoder_0/or2v0x3_1/zn 3seg_0/firseg_0/decoder_0/d4 3seg_0/firseg_0/decoder_0/or2v0x3_1/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1720 3seg_0/firseg_0/decoder_0/or2v0x3_1/a_48_39# 3seg_0/firseg_0/decoder_0/d4 3seg_0/firseg_0/decoder_0/or2v0x3_1/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1721 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_0/z 3seg_0/firseg_0/decoder_0/or2v0x3_1/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1722 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_1/zn 3seg_0/firseg_0/decoder_0/or2v0x3_1/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1723 3seg_0/firseg_0/decoder_0/or2v0x3_1/zn 3seg_0/firseg_0/decoder_0/or2v0x3_0/z gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1724 gnd 3seg_0/firseg_0/decoder_0/d4 3seg_0/firseg_0/decoder_0/or2v0x3_1/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1725 3seg_0/firseg_0/decoder_0/or2v0x3_0/z 3seg_0/firseg_0/decoder_0/or2v0x3_0/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1726 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_0/zn 3seg_0/firseg_0/decoder_0/or2v0x3_0/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1727 3seg_0/firseg_0/decoder_0/or2v0x3_0/a_31_39# 3seg_0/firseg_0/decoder_0/d0 vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1728 3seg_0/firseg_0/decoder_0/or2v0x3_0/zn 3seg_0/firseg_0/decoder_0/d2 3seg_0/firseg_0/decoder_0/or2v0x3_0/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1729 3seg_0/firseg_0/decoder_0/or2v0x3_0/a_48_39# 3seg_0/firseg_0/decoder_0/d2 3seg_0/firseg_0/decoder_0/or2v0x3_0/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1730 vdd 3seg_0/firseg_0/decoder_0/d0 3seg_0/firseg_0/decoder_0/or2v0x3_0/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1731 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_0/zn 3seg_0/firseg_0/decoder_0/or2v0x3_0/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1732 3seg_0/firseg_0/decoder_0/or2v0x3_0/zn 3seg_0/firseg_0/decoder_0/d0 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1733 gnd 3seg_0/firseg_0/decoder_0/d2 3seg_0/firseg_0/decoder_0/or2v0x3_0/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1734 decoder_0/b2 decoder_0/or2v0x3_8/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1735 vdd decoder_0/or2v0x3_8/zn decoder_0/b2 vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1736 decoder_0/or2v0x3_8/a_31_39# decoder_0/d6 vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1737 decoder_0/or2v0x3_8/zn decoder_0/or2v0x3_7/z decoder_0/or2v0x3_8/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1738 decoder_0/or2v0x3_8/a_48_39# decoder_0/or2v0x3_7/z decoder_0/or2v0x3_8/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1739 vdd decoder_0/d6 decoder_0/or2v0x3_8/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1740 gnd decoder_0/or2v0x3_8/zn decoder_0/b2 gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1741 decoder_0/or2v0x3_8/zn decoder_0/d6 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1742 gnd decoder_0/or2v0x3_7/z decoder_0/or2v0x3_8/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1743 decoder_0/or2v0x3_7/z decoder_0/or2v0x3_7/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1744 vdd decoder_0/or2v0x3_7/zn decoder_0/or2v0x3_7/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1745 decoder_0/or2v0x3_7/a_31_39# decoder_0/or2v0x3_6/z vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1746 decoder_0/or2v0x3_7/zn decoder_0/d4 decoder_0/or2v0x3_7/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1747 decoder_0/or2v0x3_7/a_48_39# decoder_0/d4 decoder_0/or2v0x3_7/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1748 vdd decoder_0/or2v0x3_6/z decoder_0/or2v0x3_7/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1749 gnd decoder_0/or2v0x3_7/zn decoder_0/or2v0x3_7/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1750 decoder_0/or2v0x3_7/zn decoder_0/or2v0x3_6/z gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1751 gnd decoder_0/d4 decoder_0/or2v0x3_7/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1752 decoder_0/or2v0x3_6/z decoder_0/or2v0x3_6/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1753 vdd decoder_0/or2v0x3_6/zn decoder_0/or2v0x3_6/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1754 decoder_0/or2v0x3_6/a_31_39# decoder_0/d3 vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1755 decoder_0/or2v0x3_6/zn decoder_0/d5 decoder_0/or2v0x3_6/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1756 decoder_0/or2v0x3_6/a_48_39# decoder_0/d5 decoder_0/or2v0x3_6/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1757 vdd decoder_0/d3 decoder_0/or2v0x3_6/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1758 gnd decoder_0/or2v0x3_6/zn decoder_0/or2v0x3_6/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1759 decoder_0/or2v0x3_6/zn decoder_0/d3 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1760 gnd decoder_0/d5 decoder_0/or2v0x3_6/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1761 decoder_0/b1 decoder_0/or2v0x3_5/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1762 vdd decoder_0/or2v0x3_5/zn decoder_0/b1 vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1763 decoder_0/or2v0x3_5/a_31_39# decoder_0/or2v0x3_4/z vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1764 decoder_0/or2v0x3_5/zn decoder_0/d6 decoder_0/or2v0x3_5/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1765 decoder_0/or2v0x3_5/a_48_39# decoder_0/d6 decoder_0/or2v0x3_5/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1766 vdd decoder_0/or2v0x3_4/z decoder_0/or2v0x3_5/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1767 gnd decoder_0/or2v0x3_5/zn decoder_0/b1 gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1768 decoder_0/or2v0x3_5/zn decoder_0/or2v0x3_4/z gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1769 gnd decoder_0/d6 decoder_0/or2v0x3_5/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1770 decoder_0/or2v0x3_4/z decoder_0/or2v0x3_4/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1771 vdd decoder_0/or2v0x3_4/zn decoder_0/or2v0x3_4/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1772 decoder_0/or2v0x3_4/a_31_39# decoder_0/d1 vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1773 decoder_0/or2v0x3_4/zn decoder_0/or2v0x3_3/z decoder_0/or2v0x3_4/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1774 decoder_0/or2v0x3_4/a_48_39# decoder_0/or2v0x3_3/z decoder_0/or2v0x3_4/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1775 vdd decoder_0/d1 decoder_0/or2v0x3_4/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1776 gnd decoder_0/or2v0x3_4/zn decoder_0/or2v0x3_4/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1777 decoder_0/or2v0x3_4/zn decoder_0/d1 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1778 gnd decoder_0/or2v0x3_3/z decoder_0/or2v0x3_4/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1779 decoder_0/or2v0x3_3/z decoder_0/or2v0x3_3/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1780 vdd decoder_0/or2v0x3_3/zn decoder_0/or2v0x3_3/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1781 decoder_0/or2v0x3_3/a_31_39# decoder_0/d5 vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1782 decoder_0/or2v0x3_3/zn decoder_0/d2 decoder_0/or2v0x3_3/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1783 decoder_0/or2v0x3_3/a_48_39# decoder_0/d2 decoder_0/or2v0x3_3/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1784 vdd decoder_0/d5 decoder_0/or2v0x3_3/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1785 gnd decoder_0/or2v0x3_3/zn decoder_0/or2v0x3_3/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1786 decoder_0/or2v0x3_3/zn decoder_0/d5 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1787 gnd decoder_0/d2 decoder_0/or2v0x3_3/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1788 decoder_0/b0 decoder_0/or2v0x3_2/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1789 vdd decoder_0/or2v0x3_2/zn decoder_0/b0 vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1790 decoder_0/or2v0x3_2/a_31_39# decoder_0/or2v0x3_1/z vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1791 decoder_0/or2v0x3_2/zn decoder_0/d6 decoder_0/or2v0x3_2/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1792 decoder_0/or2v0x3_2/a_48_39# decoder_0/d6 decoder_0/or2v0x3_2/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1793 vdd decoder_0/or2v0x3_1/z decoder_0/or2v0x3_2/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1794 gnd decoder_0/or2v0x3_2/zn decoder_0/b0 gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1795 decoder_0/or2v0x3_2/zn decoder_0/or2v0x3_1/z gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1796 gnd decoder_0/d6 decoder_0/or2v0x3_2/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1797 decoder_0/or2v0x3_1/z decoder_0/or2v0x3_1/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1798 vdd decoder_0/or2v0x3_1/zn decoder_0/or2v0x3_1/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1799 decoder_0/or2v0x3_1/a_31_39# decoder_0/or2v0x3_0/z vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1800 decoder_0/or2v0x3_1/zn decoder_0/d4 decoder_0/or2v0x3_1/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1801 decoder_0/or2v0x3_1/a_48_39# decoder_0/d4 decoder_0/or2v0x3_1/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1802 vdd decoder_0/or2v0x3_0/z decoder_0/or2v0x3_1/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1803 gnd decoder_0/or2v0x3_1/zn decoder_0/or2v0x3_1/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1804 decoder_0/or2v0x3_1/zn decoder_0/or2v0x3_0/z gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1805 gnd decoder_0/d4 decoder_0/or2v0x3_1/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
M1806 decoder_0/or2v0x3_0/z decoder_0/or2v0x3_0/zn vdd vdd pfet w=20 l=2
+ ad=160 pd=56 as=0 ps=0 
M1807 vdd decoder_0/or2v0x3_0/zn decoder_0/or2v0x3_0/z vdd pfet w=20 l=2
+ ad=0 pd=0 as=0 ps=0 
M1808 decoder_0/or2v0x3_0/a_31_39# decoder_0/d0 vdd vdd pfet w=20 l=2
+ ad=100 pd=50 as=0 ps=0 
M1809 decoder_0/or2v0x3_0/zn decoder_0/d2 decoder_0/or2v0x3_0/a_31_39# vdd pfet w=20 l=2
+ ad=148 pd=56 as=0 ps=0 
M1810 decoder_0/or2v0x3_0/a_48_39# decoder_0/d2 decoder_0/or2v0x3_0/zn vdd pfet w=16 l=2
+ ad=80 pd=42 as=0 ps=0 
M1811 vdd decoder_0/d0 decoder_0/or2v0x3_0/a_48_39# vdd pfet w=16 l=2
+ ad=0 pd=0 as=0 ps=0 
M1812 gnd decoder_0/or2v0x3_0/zn decoder_0/or2v0x3_0/z gnd nfet w=20 l=2
+ ad=0 pd=0 as=126 ps=54 
M1813 decoder_0/or2v0x3_0/zn decoder_0/d0 gnd gnd nfet w=10 l=2
+ ad=80 pd=36 as=0 ps=0 
M1814 gnd decoder_0/d2 decoder_0/or2v0x3_0/zn gnd nfet w=10 l=2
+ ad=0 pd=0 as=0 ps=0 
C0 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z 30.2fF
C1 3seg_0/firseg_0/comp_0/an2v0x2_1/b 3seg_0/firseg_0/decoder_0/b0 2.2fF
C2 3seg_0/2seg_0/an2v0x3_0/z 3seg_0/2seg_0/1counter_0/or2v0x3_1/a 2.1fF
C3 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/bn 9.1fF
C4 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/sn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# 9.2fF
C5 decoder_0/b2 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/zn 2.7fF
C6 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# 3seg_0/firseg_0/decoder_0/b2 4.8fF
C7 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/zn vdd 12.7fF
C8 gnd 3seg_0/2seg_0/or3v0x3_0/zn 12.2fF
C9 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/zn 9.3fF
C10 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# 3seg_0/2seg_0/or3v0x3_0/b 5.0fF
C11 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/sn 9.2fF
C12 vdd 3seg_0/2seg_0/iv1v0x3_0/a 15.3fF
C13 3seg_0/2seg_0/ud 3seg_0/2seg_0/1counter_0/an2v0x3_0/zn 2.6fF
C14 decoder_0/or2v0x3_1/z decoder_0/or2v0x3_0/z 4.6fF
C15 gnd 3seg_0/firseg_0/comp_0/an2v0x2_4/zn 8.9fF
C16 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/zn 2.2fF
C17 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an 3.3fF
C18 3seg_0/2seg_0/totdiff3_0/mux_0/b1 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# 6.6fF
C19 gnd 3seg_0/firseg_0/decoder_0/d4 68.9fF
C20 3seg_0/firseg_0/comp_0/an3v0x2_0/zn gnd 8.8fF
C21 vdd 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/bn 13.7fF
C22 gnd decoder_0/or2v0x3_7/zn 9.0fF
C23 3seg_0/2seg_0/totdiff3_0/mux_0/b1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn 2.7fF
C24 gnd 3seg_0/firseg_0/decoder_0/d2 23.3fF
C25 3seg_0/2seg_0/an2v0x3_0/b vdd 6.5fF
C26 gnd 3seg_0/2seg_0/ud 27.9fF
C27 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/sn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# 9.3fF
C28 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/bn 9.1fF
C29 decoder_0/or2v0x3_4/zn vdd 12.7fF
C30 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_2/b 23.4fF
C31 gnd 3seg_0/firseg_0/comp_0/an2v0x2_2/zn 8.9fF
C32 gnd decoder_0/b1 15.9fF
C33 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/an 9.5fF
C34 gnd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/cn 17.1fF
C35 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_1/zn 9.5fF
C36 gnd decoder_0/d4 68.9fF
C37 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn 4.5fF
C38 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 11.9fF
C39 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/iz 24.9fF
C40 gnd 3seg_0/firseg_0/comp_0/nd3v0x2_0/c 18.9fF
C41 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn 18.9fF
C42 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/zn 9.3fF
C43 3seg_0/2seg_0/totdiff3_0/mux_0/b1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an 3.9fF
C44 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn 4.5fF
C45 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z 34.4fF
C46 vdd 3seg_0/firseg_0/decoder_0/d3 28.2fF
C47 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z 3seg_0/2seg_0/1counter_0/bf1v0x4_0/w_n4_n4# 2.0fF
C48 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_1/zn 9.0fF
C49 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/zn 8.9fF
C50 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/zn 8.9fF
C51 3seg_0/2seg_0/an2v0x3_0/z 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/an 2.6fF
C52 3seg_0/firseg_0/decoder_0/b0 3seg_0/firseg_0/decoder_0/or2v0x3_1/z 4.7fF
C53 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/bn 3seg_0/firseg_0/3_bitmux_0/o2 2.6fF
C54 gnd decoder_0/b0 10.9fF
C55 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/zn 4.4fF
C56 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/zn 9.3fF
C57 3seg_0/firseg_0/out 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# 18.7fF
C58 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a 12.4fF
C59 gnd 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/d 13.6fF
C60 vdd 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/bn 13.7fF
C61 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn vdd 18.9fF
C62 gnd decoder_0/d6 48.5fF
C63 gnd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n1 9.9fF
C64 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/z 12.8fF
C65 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/zn 8.9fF
C66 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 3seg_0/firseg_0/comp_0/nr3v0x2_0/a 15.0fF
C67 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_3/b 15.2fF
C68 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_2/zn 13.3fF
C69 3seg_0/2seg_0/totdiff3_0/mux_0/b2 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn 2.7fF
C70 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/in_2c 34.0fF
C71 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/b0 26.2fF
C72 gnd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/d 13.6fF
C73 gnd 3seg_0/firseg_0/decoder_0/b2 37.2fF
C74 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_1/w_n4_n4# 19.0fF
C75 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/in_2c 17.8fF
C76 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/sn 9.3fF
C77 decoder_0/or2v0x3_1/z decoder_0/or2v0x3_2/zn 2.0fF
C78 vdd decoder_0/or2v0x3_7/z 11.4fF
C79 3seg_0/firseg_0/decoder_0/or2v0x3_2/zn 3seg_0/firseg_0/decoder_0/b0 2.2fF
C80 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/zn 8.9fF
C81 3seg_0/2seg_0/1counter_0/an2v0x3_0/zn vdd 13.3fF
C82 3seg_0/firseg_0/decoder_0/or2v0x3_6/z gnd 9.2fF
C83 3seg_0/firseg_0/decoder_0/b0 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# 11.6fF
C84 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn 18.8fF
C85 gnd 3seg_0/firseg_0/comp_0/an2v0x2_0/b 32.8fF
C86 3seg_0/firseg_0/comp_0/an3v0x2_0/zn 3seg_0/firseg_0/comp_0/an3v0x2_1/a 2.5fF
C87 3seg_0/2seg_0/or3v0x3_0/a 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# 5.2fF
C88 3seg_0/2seg_0/an2v0x3_0/a vdd 8.1fF
C89 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 3seg_0/firseg_0/out 5.6fF
C90 3seg_0/firseg_0/out 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# 30.3fF
C91 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/z 10.2fF
C92 gnd 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/an 9.2fF
C93 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn 19.1fF
C94 3seg_0/firseg_0/decoder_0/or2v0x3_2/zn 3seg_0/firseg_0/decoder_0/or2v0x3_1/z 2.0fF
C95 3seg_0/firseg_0/decoder_0/or2v0x3_0/zn 3seg_0/firseg_0/decoder_0/or2v0x3_0/z 2.3fF
C96 gnd vdd 48.3fF
C97 gnd 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/ci 27.5fF
C98 gnd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/cn 17.1fF
C99 gnd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n4 7.3fF
C100 vdd decoder_0/or2v0x3_6/zn 12.7fF
C101 3seg_0/firseg_0/out 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# 36.4fF
C102 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/zn 3seg_0/2seg_0/totdiff3_0/mux_0/b2 2.7fF
C103 vdd 3seg_0/firseg_0/comp_0/an2v0x2_4/z 10.7fF
C104 gnd 3seg_0/2seg_0/1counter_0/or2v0x3_1/zn 9.0fF
C105 vdd decoder_0/or2v0x3_5/zn 12.7fF
C106 3seg_0/firseg_0/decoder_0/or2v0x3_4/zn 3seg_0/firseg_0/decoder_0/d6 2.1fF
C107 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/bn 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/d 2.8fF
C108 gnd decoder_0/d5 20.2fF
C109 gnd decoder_0/or2v0x3_6/z 9.2fF
C110 vdd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/ci 16.6fF
C111 3seg_0/firseg_0/decoder_0/or2v0x3_7/z vdd 11.4fF
C112 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an 25.5fF
C113 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/zn 8.8fF
C114 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn 4.5fF
C115 gnd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n4 7.3fF
C116 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n1 vdd 8.4fF
C117 gnd decoder_0/d1 7.6fF
C118 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 3seg_0/firseg_0/decoder_0/b0 8.1fF
C119 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 3seg_0/firseg_0/comp_0/an3v0x2_1/zn 5.8fF
C120 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a gnd 20.0fF
C121 3seg_0/firseg_0/decoder_0/b0 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# 4.8fF
C122 vdd 3seg_0/2seg_0/1counter_0/or2v0x3_0/zn 12.7fF
C123 decoder_0/b2 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# 8.7fF
C124 3seg_0/firseg_0/comp_0/an3v0x2_2/b 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 21.4fF
C125 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn 18.7fF
C126 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/an vdd 9.9fF
C127 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/mux_0/a0 4.1fF
C128 gnd decoder_0/or2v0x3_1/zn 9.0fF
C129 gnd decoder_0/or2v0x3_3/z 12.6fF
C130 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/zn 8.9fF
C131 3seg_0/2seg_0/an2v0x3_0/z 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/ci 2.2fF
C132 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/a0 35.2fF
C133 vdd decoder_0/d0 14.1fF
C134 gnd 3seg_0/firseg_0/comp_0/an3v0x2_0/z 36.9fF
C135 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/mux_0/a2 4.6fF
C136 gnd 3seg_0/firseg_0/comp_0/an2v0x2_3/z 20.8fF
C137 gnd 3seg_0/firseg_0/comp_0/an3v0x2_2/zn 8.8fF
C138 vdd 3seg_0/2seg_0/or3v0x3_0/b 8.0fF
C139 gnd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/d 13.6fF
C140 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/bn 6.7fF
C141 3seg_0/firseg_0/comp_0/an3v0x2_1/a 3seg_0/firseg_0/comp_0/an2v0x2_0/b 2.5fF
C142 3seg_0/2seg_0/totdiff3_0/mux_0/b1 vdd 13.1fF
C143 gnd 3seg_0/firseg_0/comp_0/an3v0x2_3/zn 8.8fF
C144 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/an 9.5fF
C145 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# 2.3fF
C146 vdd 3seg_0/firseg_0/decoder_0/d1 17.9fF
C147 vdd 3seg_0/2seg_0/1counter_0/or2v0x3_1/a 23.6fF
C148 3seg_0/firseg_0/decoder_0/or2v0x3_6/z 3seg_0/firseg_0/decoder_0/or2v0x3_7/zn 2.0fF
C149 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 3seg_0/firseg_0/comp_0/nr3v0x2_0/z 21.8fF
C150 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/a 40.8fF
C151 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n2 vdd 12.4fF
C152 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/zn 8.9fF
C153 vdd 3seg_0/firseg_0/comp_0/an3v0x2_1/a 72.4fF
C154 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# 5.0fF
C155 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/zn 4.4fF
C156 gnd decoder_0/or2v0x3_3/zn 9.0fF
C157 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn 11.2fF
C158 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_7/zn 12.7fF
C159 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_3/zn 9.5fF
C160 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn 31.6fF
C161 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/b 20.5fF
C162 vdd 3seg_0/firseg_0/comp_0/an2v0x2_2/z 9.4fF
C163 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a 25.9fF
C164 gnd 3seg_0/firseg_0/decoder_0/d5 20.2fF
C165 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/a2 14.9fF
C166 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/firseg_0/decoder_0/b0 2.3fF
C167 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a 2.1fF
C168 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 3seg_0/firseg_0/comp_0/nd3v0x2_0/a 6.2fF
C169 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# 3seg_0/firseg_0/3_bitmux_0/o2 6.3fF
C170 3seg_0/firseg_0/decoder_0/or2v0x3_1/z 3seg_0/firseg_0/decoder_0/or2v0x3_0/z 4.6fF
C171 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn 3.3fF
C172 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n4 gnd 7.3fF
C173 gnd decoder_0/b2 11.2fF
C174 3seg_0/firseg_0/comp_0/or3v0x2_0/zn vdd 9.0fF
C175 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/zn vdd 8.8fF
C176 3seg_0/2seg_0/or3v0x3_0/a_57_38# 3seg_0/2seg_0/or3v0x3_0/a 2.6fF
C177 3seg_0/firseg_0/decoder_0/b1 3seg_0/firseg_0/decoder_0/d6 2.7fF
C178 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# 3seg_0/firseg_0/decoder_0/b1 4.8fF
C179 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/iz 25.5fF
C180 gnd 3seg_0/2seg_0/1counter_0/or2v0x3_0/z 9.7fF
C181 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_3/zn 9.0fF
C182 vdd 3seg_0/firseg_0/comp_0/an2v0x2_1/z 22.0fF
C183 gnd 3seg_0/2seg_0/or3v0x3_0/c 6.7fF
C184 vdd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n2 12.4fF
C185 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# 3seg_0/firseg_0/decoder_0/b1 13.4fF
C186 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/z vdd 2.4fF
C187 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/z 24.6fF
C188 gnd 3seg_0/2seg_0/1counter_0/or2v0x3_1/z 10.5fF
C189 3seg_0/2seg_0/ud 3seg_0/2seg_0/iv1v0x3_0/z 3.1fF
C190 vdd 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/an 6.0fF
C191 decoder_0/b0 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/zn 2.7fF
C192 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a 59.6fF
C193 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/b2 11.9fF
C194 gnd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n2 7.2fF
C195 3seg_0/firseg_0/comp_0/an3v0x2_0/zn 3seg_0/firseg_0/decoder_0/b0 4.6fF
C196 3seg_0/firseg_0/comp_0/nr3v0x2_0/a 3seg_0/firseg_0/decoder_0/b2 2.5fF
C197 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/cn vdd 46.5fF
C198 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_0/zn 12.7fF
C199 3seg_0/firseg_0/out decoder_0/b0 3.2fF
C200 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z 3seg_0/2seg_0/1counter_0/bf1v0x4_2/w_n4_n4# 2.0fF
C201 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/zn vdd 10.2fF
C202 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z 29.8fF
C203 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a 3seg_0/firseg_0/3_bitmux_0/o0 2.0fF
C204 3seg_0/2seg_0/ud 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# 18.7fF
C205 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# 3seg_0/2seg_0/totdiff3_0/mux_0/a1 13.4fF
C206 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/or2v0x3_0/zn 9.0fF
C207 vdd decoder_0/or2v0x3_0/z 19.2fF
C208 3seg_0/2seg_0/totdiff3_0/mux_0/b2 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an 3.9fF
C209 3seg_0/2seg_0/totdiff3_0/mux_0/b0 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# 8.7fF
C210 3seg_0/2seg_0/ud 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# 15.6fF
C211 gnd 3seg_0/2seg_0/iv1v0x3_0/a 7.6fF
C212 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# 5.2fF
C213 3seg_0/firseg_0/decoder_0/b0 decoder_0/b1 2.9fF
C214 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/bn 2.6fF
C215 vdd 3seg_0/firseg_0/comp_0/nr3v0x2_0/a 4.0fF
C216 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/b 20.5fF
C217 gnd 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/bn 6.5fF
C218 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/z 24.6fF
C219 gnd 3seg_0/2seg_0/an2v0x3_0/b 5.5fF
C220 vdd 3seg_0/firseg_0/comp_0/or3v0x2_1/zn 9.0fF
C221 vdd decoder_0/or2v0x3_0/zn 12.7fF
C222 decoder_0/b0 decoder_0/or2v0x3_2/zn 2.2fF
C223 3seg_0/firseg_0/decoder_0/or2v0x3_5/zn vdd 12.7fF
C224 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c 40.7fF
C225 gnd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# 25.5fF
C226 decoder_0/or2v0x3_4/zn gnd 9.0fF
C227 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c vdd 39.6fF
C228 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/zn 12.7fF
C229 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/bn 15.4fF
C230 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/zn 2.2fF
C231 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_2/b 21.8fF
C232 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# 76.0fF
C233 3seg_0/firseg_0/decoder_0/or2v0x3_3/zn 3seg_0/firseg_0/decoder_0/d1 3.7fF
C234 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/b vdd 20.5fF
C235 vdd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n1 8.4fF
C236 decoder_0/or2v0x3_1/zn decoder_0/or2v0x3_0/z 2.0fF
C237 3seg_0/2seg_0/1counter_0/bf1v0x4_0/w_n4_n4# 3seg_0/2seg_0/1counter_0/bf1v0x4_0/an 9.7fF
C238 3seg_0/firseg_0/decoder_0/or2v0x3_1/z 3seg_0/firseg_0/decoder_0/or2v0x3_1/zn 2.3fF
C239 3seg_0/2seg_0/1counter_0/bf1v0x4_1/w_n4_n4# 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a 3.9fF
C240 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/sn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# 9.3fF
C241 3seg_0/firseg_0/comp_0/an2v0x2_1/b vdd 14.2fF
C242 3seg_0/firseg_0/out vdd 10.6fF
C243 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn 13.9fF
C244 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/iz vdd 15.8fF
C245 3seg_0/firseg_0/comp_0/nr2v0x2_1/a 3seg_0/firseg_0/comp_0/nd3v0x2_0/c 3.8fF
C246 gnd 3seg_0/firseg_0/decoder_0/d3 7.6fF
C247 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/an 9.9fF
C248 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# 2.3fF
C249 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 4.3fF
C250 decoder_0/d2 vdd 16.1fF
C251 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/zn 11.9fF
C252 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 3seg_0/firseg_0/comp_0/an3v0x2_2/z 21.1fF
C253 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a 20.0fF
C254 3seg_0/2seg_0/1counter_0/an2v0x3_1/b vdd 20.2fF
C255 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/z vdd 17.9fF
C256 gnd 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/bn 6.5fF
C257 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_4/zn 12.7fF
C258 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn 11.9fF
C259 vdd 3seg_0/2seg_0/iv1v0x3_0/z 5.9fF
C260 3seg_0/firseg_0/decoder_0/b0 3seg_0/firseg_0/comp_0/an2v0x2_0/b 4.9fF
C261 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_2/zn 9.5fF
C262 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a 2.1fF
C263 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a 37.1fF
C264 3seg_0/firseg_0/comp_0/nr3v0x2_0/a 3seg_0/firseg_0/comp_0/an3v0x2_2/zn 2.1fF
C265 3seg_0/firseg_0/decoder_0/d0 3seg_0/firseg_0/decoder_0/or2v0x3_0/z 3.9fF
C266 3seg_0/firseg_0/comp_0/an3v0x2_2/b 3seg_0/firseg_0/comp_0/an2v0x2_0/b 2.5fF
C267 vdd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/ci 16.6fF
C268 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/b0 10.9fF
C269 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/bn 14.4fF
C270 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/in_2c 17.5fF
C271 3seg_0/2seg_0/totdiff3_0/mux_0/a0 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# 4.8fF
C272 decoder_0/or2v0x3_1/z decoder_0/b0 4.7fF
C273 vdd decoder_0/or2v0x3_2/zn 12.7fF
C274 vdd 3seg_0/firseg_0/decoder_0/b0 47.8fF
C275 vdd 3seg_0/firseg_0/comp_0/an3v0x2_1/zn 4.9fF
C276 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# 20.7fF
C277 3seg_0/2seg_0/totdiff3_0/mux_0/a0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn 4.6fF
C278 vdd 3seg_0/firseg_0/comp_0/an2v0x2_1/zn 8.8fF
C279 3seg_0/firseg_0/comp_0/an3v0x2_2/b vdd 39.7fF
C280 decoder_0/b0 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# 6.6fF
C281 gnd decoder_0/or2v0x3_7/z 15.6fF
C282 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 3seg_0/2seg_0/totdiff3_0/mux_0/a1 4.6fF
C283 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_0/zn 9.5fF
C284 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/zn 8.8fF
C285 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/zn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# 8.9fF
C286 3seg_0/2seg_0/or3v0x3_0/b 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# 2.3fF
C287 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an 3.3fF
C288 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/bn 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/d 2.8fF
C289 vdd decoder_0/or2v0x3_4/z 18.3fF
C290 vdd decoder_0/or2v0x3_8/zn 12.7fF
C291 gnd 3seg_0/2seg_0/an2v0x3_0/a 11.5fF
C292 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_1/z 19.4fF
C293 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/sn 3seg_0/2seg_0/or3v0x3_0/a 4.3fF
C294 3seg_0/2seg_0/totdiff3_0/mux_0/b1 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# 10.2fF
C295 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/w_n4_n4# 18.2fF
C296 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/zn 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z 2.2fF
C297 3seg_0/2seg_0/totdiff3_0/mux_0/b0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn 2.7fF
C298 vdd 3seg_0/firseg_0/comp_0/nr2v0x2_1/a 7.1fF
C299 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/w_n4_n4# 18.8fF
C300 gnd decoder_0/or2v0x3_6/zn 9.0fF
C301 decoder_0/b1 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# 10.2fF
C302 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/bn 14.4fF
C303 3seg_0/firseg_0/decoder_0/or2v0x3_6/zn vdd 12.7fF
C304 gnd 3seg_0/firseg_0/comp_0/an2v0x2_4/z 9.8fF
C305 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 3seg_0/firseg_0/comp_0/nd3v0x2_0/c 5.7fF
C306 gnd decoder_0/or2v0x3_5/zn 9.0fF
C307 3seg_0/firseg_0/3_bitmux_0/o1 vdd 53.3fF
C308 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# decoder_0/b1 6.6fF
C309 gnd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/ci 27.5fF
C310 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/z 17.9fF
C311 3seg_0/firseg_0/decoder_0/or2v0x3_7/z gnd 15.6fF
C312 decoder_0/b0 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# 8.7fF
C313 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a vdd 12.4fF
C314 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/an 21.6fF
C315 vdd 3seg_0/firseg_0/comp_0/nr3v0x2_0/z 8.7fF
C316 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/zn 8.9fF
C317 decoder_0/or2v0x3_1/z vdd 19.4fF
C318 gnd 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n1 9.9fF
C319 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_2/zn 12.7fF
C320 gnd 3seg_0/2seg_0/1counter_0/or2v0x3_0/zn 9.0fF
C321 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# 3seg_0/2seg_0/ud 36.4fF
C322 vdd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# 20.7fF
C323 vdd 3seg_0/2seg_0/or3v0x3_0/a 15.7fF
C324 3seg_0/2seg_0/totdiff3_0/mux_0/b1 3seg_0/2seg_0/totdiff3_0/mux_0/b0 18.4fF
C325 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/bn 11.2fF
C326 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/an 5.5fF
C327 vdd 3seg_0/firseg_0/3_bitmux_0/o2 53.4fF
C328 vdd 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/bn 13.7fF
C329 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/a0 14.9fF
C330 3seg_0/firseg_0/decoder_0/or2v0x3_0/z 3seg_0/firseg_0/decoder_0/d2 2.2fF
C331 gnd decoder_0/d0 7.6fF
C332 vdd 3seg_0/firseg_0/comp_0/an2v0x2_3/b 13.7fF
C333 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 3seg_0/firseg_0/decoder_0/b2 11.6fF
C334 vdd 3seg_0/firseg_0/comp_0/nd3v0x2_0/a 9.6fF
C335 3seg_0/2seg_0/ud 3seg_0/2seg_0/an2v0x3_0/zn 2.7fF
C336 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/a1 38.6fF
C337 vdd 3seg_0/firseg_0/comp_0/an2v0x2_0/zn 8.8fF
C338 vdd decoder_0/d3 30.9fF
C339 gnd 3seg_0/2seg_0/or3v0x3_0/b 16.8fF
C340 vdd 3seg_0/firseg_0/decoder_0/b1 55.2fF
C341 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# 3seg_0/firseg_0/decoder_0/b2 11.6fF
C342 decoder_0/or2v0x3_1/z decoder_0/or2v0x3_1/zn 2.3fF
C343 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/a 34.7fF
C344 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/sn 9.3fF
C345 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a 3seg_0/firseg_0/3_bitmux_0/o2 2.0fF
C346 3seg_0/2seg_0/1counter_0/bf1v0x4_2/an 3seg_0/2seg_0/1counter_0/bf1v0x4_2/w_n4_n4# 9.7fF
C347 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/bn 2.6fF
C348 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/sn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_32# 9.3fF
C349 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/b1 17.2fF
C350 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/sn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# 9.2fF
C351 vdd 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/a 6.0fF
C352 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_2/a 15.5fF
C353 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_4/z 18.3fF
C354 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# vdd 87.6fF
C355 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_3/z 12.1fF
C356 vdd 3seg_0/firseg_0/decoder_0/d6 35.0fF
C357 gnd 3seg_0/firseg_0/decoder_0/d1 7.6fF
C358 gnd 3seg_0/2seg_0/1counter_0/or2v0x3_1/a 9.3fF
C359 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/a 18.1fF
C360 3seg_0/2seg_0/1counter_0/bf1v0x4_0/w_n4_n4# 3seg_0/2seg_0/1counter_0/bf1v0x4_0/a 3.9fF
C361 3seg_0/firseg_0/decoder_0/or2v0x3_0/z 3seg_0/firseg_0/decoder_0/or2v0x3_1/zn 2.0fF
C362 gnd 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n2 7.2fF
C363 gnd 3seg_0/firseg_0/comp_0/an3v0x2_1/a 57.3fF
C364 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# 3seg_0/2seg_0/totdiff3_0/mux_0/a2 4.8fF
C365 vdd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# 59.4fF
C366 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/zn 11.9fF
C367 3seg_0/2seg_0/an2v0x3_0/z vdd 59.1fF
C368 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_7/zn 9.0fF
C369 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/zn 8.8fF
C370 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_8/zn 12.7fF
C371 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/an 9.9fF
C372 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn 18.8fF
C373 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/b 5.9fF
C374 gnd 3seg_0/firseg_0/comp_0/an2v0x2_2/z 11.1fF
C375 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a 2.3fF
C376 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/bn 2.4fF
C377 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# 3seg_0/2seg_0/or3v0x3_0/c 2.3fF
C378 3seg_0/firseg_0/decoder_0/d0 vdd 14.1fF
C379 3seg_0/firseg_0/comp_0/an2v0x2_3/zn vdd 8.8fF
C380 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/sn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# 9.2fF
C381 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/zn vdd 4.4fF
C382 gnd 3seg_0/firseg_0/comp_0/or3v0x2_0/zn 10.9fF
C383 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/zn 8.9fF
C384 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a 59.6fF
C385 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/zn 8.9fF
C386 3seg_0/firseg_0/out 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# 15.2fF
C387 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# vdd 59.4fF
C388 gnd 3seg_0/firseg_0/comp_0/an2v0x2_1/z 8.7fF
C389 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/zn vdd 12.7fF
C390 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/zn 10.3fF
C391 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn 17.7fF
C392 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# 3seg_0/2seg_0/totdiff3_0/mux_0/b2 8.7fF
C393 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 3seg_0/firseg_0/comp_0/an3v0x2_0/z 9.5fF
C394 vdd 3seg_0/firseg_0/comp_0/an3v0x2_3/z 15.4fF
C395 vdd 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/an 6.0fF
C396 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_1/a 15.5fF
C397 gnd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n2 7.2fF
C398 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/zn 9.3fF
C399 3seg_0/firseg_0/comp_0/an3v0x2_3/zn 3seg_0/firseg_0/decoder_0/b1 3.6fF
C400 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/z 2.5fF
C401 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/z 12.8fF
C402 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 3seg_0/firseg_0/comp_0/an3v0x2_2/zn 5.8fF
C403 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/zn 3.1fF
C404 gnd 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/an 9.2fF
C405 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z 3seg_0/2seg_0/1counter_0/bf1v0x4_1/w_n4_n4# 3.3fF
C406 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a 25.9fF
C407 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_0/z 19.2fF
C408 vdd 3seg_0/2seg_0/an2v0x3_0/zn 13.3fF
C409 gnd 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/cn 17.1fF
C410 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_0/zn 9.0fF
C411 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_2/z 12.7fF
C412 gnd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/zn 20.1fF
C413 vdd 3seg_0/firseg_0/3_bitmux_0/o0 53.4fF
C414 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an 25.5fF
C415 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an 27.4fF
C416 3seg_0/2seg_0/an2v0x3_0/z 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/d 2.4fF
C417 3seg_0/2seg_0/ud 3seg_0/2seg_0/1counter_0/an2v0x3_3/b 2.4fF
C418 vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/z 3.3fF
C419 gnd decoder_0/or2v0x3_0/z 10.3fF
C420 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z vdd 35.1fF
C421 decoder_0/d6 decoder_0/b1 2.7fF
C422 gnd 3seg_0/firseg_0/comp_0/nr3v0x2_0/a 19.9fF
C423 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/b 7.3fF
C424 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/bn 15.4fF
C425 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/z 12.8fF
C426 3seg_0/2seg_0/or3v0x3_0/zn vdd 13.4fF
C427 gnd 3seg_0/firseg_0/comp_0/or3v0x2_1/zn 10.9fF
C428 gnd decoder_0/or2v0x3_0/zn 9.0fF
C429 3seg_0/firseg_0/decoder_0/or2v0x3_5/zn gnd 9.0fF
C430 vdd 3seg_0/firseg_0/comp_0/an2v0x2_4/zn 8.8fF
C431 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c 35.0fF
C432 3seg_0/2seg_0/1counter_0/an2v0x3_3/b 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z 2.9fF
C433 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/zn 8.9fF
C434 3seg_0/firseg_0/comp_0/an3v0x2_0/zn vdd 10.7fF
C435 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c gnd 34.1fF
C436 vdd 3seg_0/firseg_0/decoder_0/d4 15.8fF
C437 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/sn 3seg_0/firseg_0/3_bitmux_0/o0 4.3fF
C438 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/or2v0x3_0/zn 9.0fF
C439 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/bn 9.1fF
C440 vdd decoder_0/or2v0x3_7/zn 12.7fF
C441 vdd 3seg_0/firseg_0/decoder_0/d2 16.1fF
C442 3seg_0/firseg_0/decoder_0/or2v0x3_3/zn 3seg_0/firseg_0/decoder_0/d6 2.2fF
C443 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/b 5.9fF
C444 gnd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n1 9.9fF
C445 3seg_0/firseg_0/comp_0/or3v0x2_0/zn 3seg_0/firseg_0/comp_0/an3v0x2_1/a 4.1fF
C446 3seg_0/2seg_0/ud vdd 30.0fF
C447 gnd 3seg_0/firseg_0/comp_0/an2v0x2_1/b 5.9fF
C448 gnd 3seg_0/firseg_0/out 14.6fF
C449 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/iz gnd 24.9fF
C450 decoder_0/b2 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# 6.6fF
C451 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/bn 15.4fF
C452 decoder_0/d0 decoder_0/or2v0x3_0/z 3.9fF
C453 decoder_0/or2v0x3_6/z decoder_0/or2v0x3_7/zn 2.0fF
C454 3seg_0/2seg_0/totdiff3_0/mux_0/b0 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# 6.6fF
C455 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n4 3seg_0/2seg_0/an2v0x3_0/z 2.3fF
C456 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/an 5.5fF
C457 decoder_0/d2 gnd 23.3fF
C458 3seg_0/2seg_0/an2v0x3_0/z 3seg_0/2seg_0/1counter_0/or2v0x3_0/z 2.7fF
C459 vdd 3seg_0/firseg_0/comp_0/an2v0x2_2/zn 8.8fF
C460 vdd decoder_0/b1 14.6fF
C461 vdd 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/cn 46.5fF
C462 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_1/zn 13.3fF
C463 vdd decoder_0/d4 17.1fF
C464 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/zn 18.9fF
C465 3seg_0/2seg_0/1counter_0/bf1v0x4_1/w_n4_n4# 3seg_0/2seg_0/1counter_0/bf1v0x4_1/an 9.7fF
C466 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/iz 15.8fF
C467 vdd 3seg_0/firseg_0/comp_0/nd3v0x2_0/c 5.0fF
C468 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_1/b 10.0fF
C469 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/z 10.2fF
C470 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_4/zn 9.0fF
C471 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# 3seg_0/2seg_0/totdiff3_0/mux_0/a2 11.6fF
C472 gnd 3seg_0/2seg_0/iv1v0x3_0/z 4.5fF
C473 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_2/w_n4_n4# 3seg_0/firseg_0/3_bitmux_0/o2 2.3fF
C474 3seg_0/2seg_0/totdiff3_0/mux_0/b0 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/zn 2.7fF
C475 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z 39.1fF
C476 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_1/zn 12.7fF
C477 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/zn 8.8fF
C478 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/zn 8.8fF
C479 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a 18.1fF
C480 3seg_0/2seg_0/or3v0x3_0/a 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# 2.3fF
C481 3seg_0/firseg_0/3_bitmux_0/o1 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/a 2.0fF
C482 vdd decoder_0/b0 16.6fF
C483 gnd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/ci 27.5fF
C484 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn 2.3fF
C485 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xnr2v8x05_0/bn 6.7fF
C486 vdd 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/d 9.8fF
C487 gnd decoder_0/or2v0x3_2/zn 9.0fF
C488 gnd 3seg_0/firseg_0/decoder_0/b0 64.1fF
C489 vdd decoder_0/d6 35.0fF
C490 gnd 3seg_0/firseg_0/comp_0/an3v0x2_1/zn 8.8fF
C491 vdd 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/z 24.6fF
C492 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# 3seg_0/2seg_0/or3v0x3_0/c 6.3fF
C493 vdd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n1 8.4fF
C494 gnd 3seg_0/firseg_0/comp_0/an2v0x2_1/zn 8.9fF
C495 vdd 3seg_0/2seg_0/1counter_0/an2v0x3_3/b 34.2fF
C496 gnd 3seg_0/firseg_0/comp_0/an3v0x2_2/b 23.0fF
C497 vdd 3seg_0/2seg_0/1counter_0/bf1v0x4_1/an 9.5fF
C498 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# 3seg_0/2seg_0/totdiff3_0/mux_0/a1 4.8fF
C499 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# 25.3fF
C500 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/zn 9.3fF
C501 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/zn 10.8fF
C502 gnd decoder_0/or2v0x3_4/z 9.2fF
C503 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/d vdd 9.8fF
C504 gnd decoder_0/or2v0x3_8/zn 9.0fF
C505 vdd 3seg_0/firseg_0/decoder_0/b2 31.1fF
C506 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_1/w_n4_32# 3seg_0/2seg_0/totdiff3_0/mux_0/b2 6.6fF
C507 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_1/z 10.3fF
C508 3seg_0/2seg_0/totdiff3_0/diff2_2/in_2c vdd 33.2fF
C509 3seg_0/2seg_0/1counter_0/or2v0x3_1/z 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/an 3.7fF
C510 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/zn 3seg_0/firseg_0/3_bitmux_0/o2 4.3fF
C511 3seg_0/2seg_0/an2v0x3_0/z 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/bn 4.7fF
C512 3seg_0/firseg_0/decoder_0/or2v0x3_6/z vdd 20.6fF
C513 gnd 3seg_0/firseg_0/comp_0/nr2v0x2_1/a 22.9fF
C514 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/zn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# 8.9fF
C515 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn vdd 31.6fF
C516 vdd 3seg_0/firseg_0/comp_0/an2v0x2_0/b 49.9fF
C517 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/bn 7.5fF
C518 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/zn 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c 3.1fF
C519 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_6/zn 9.0fF
C520 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/sn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# 9.2fF
C521 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/z vdd 17.9fF
C522 3seg_0/2seg_0/totdiff3_0/mux_0/a0 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_32# 11.6fF
C523 vdd 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/an 6.0fF
C524 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn 31.6fF
C525 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/zn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# 9.3fF
C526 3seg_0/firseg_0/3_bitmux_0/o1 gnd 60.5fF
C527 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/ci vdd 16.6fF
C528 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/z 10.2fF
C529 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/cn vdd 46.5fF
C530 vdd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n4 8.9fF
C531 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/a 20.0fF
C532 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/sn 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_1/w_n4_32# 9.3fF
C533 gnd 3seg_0/firseg_0/comp_0/nr3v0x2_0/z 21.2fF
C534 decoder_0/or2v0x3_1/z gnd 10.3fF
C535 vdd 3seg_0/2seg_0/1counter_0/or2v0x3_1/zn 12.7fF
C536 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_2/zn 9.0fF
C537 vdd decoder_0/d5 23.0fF
C538 decoder_0/or2v0x3_6/z vdd 20.6fF
C539 3seg_0/2seg_0/ud 3seg_0/2seg_0/totdiff3_0/mux_0/a2 4.5fF
C540 gnd 3seg_0/2seg_0/or3v0x3_0/a 8.1fF
C541 gnd 3seg_0/2seg_0/1counter_0/tf_1/xor2v0x05_0/bn 6.5fF
C542 gnd 3seg_0/firseg_0/3_bitmux_0/o2 60.5fF
C543 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/ci 3seg_0/2seg_0/1counter_0/bf1v0x4_0/a 2.1fF
C544 vdd decoder_0/d1 17.9fF
C545 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/n4 vdd 8.9fF
C546 gnd 3seg_0/firseg_0/comp_0/an2v0x2_3/b 15.0fF
C547 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/a vdd 12.4fF
C548 gnd 3seg_0/firseg_0/comp_0/nd3v0x2_0/a 21.8fF
C549 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/bn 2.4fF
C550 3seg_0/firseg_0/decoder_0/b0 3seg_0/firseg_0/comp_0/an3v0x2_1/a 6.8fF
C551 gnd 3seg_0/2seg_0/totdiff3_0/mux_0/a1 15.3fF
C552 vdd decoder_0/or2v0x3_1/zn 12.7fF
C553 vdd decoder_0/or2v0x3_3/z 12.1fF
C554 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_1/zn 8.8fF
C555 gnd 3seg_0/firseg_0/comp_0/an2v0x2_0/zn 8.9fF
C556 gnd decoder_0/d3 7.6fF
C557 gnd 3seg_0/firseg_0/decoder_0/b1 21.2fF
C558 3seg_0/2seg_0/1counter_0/bf1v0x4_2/a 3seg_0/2seg_0/1counter_0/bf1v0x4_2/w_n4_n4# 3.9fF
C559 3seg_0/firseg_0/comp_0/an3v0x2_2/b 3seg_0/firseg_0/comp_0/an3v0x2_1/a 5.2fF
C560 decoder_0/or2v0x3_3/zn decoder_0/d6 2.2fF
C561 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/sn 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_2/w_n4_n4# 9.2fF
C562 vdd 3seg_0/firseg_0/comp_0/an3v0x2_0/z 2.3fF
C563 gnd 3seg_0/2seg_0/1counter_0/bf1v0x4_2/a 18.1fF
C564 3seg_0/2seg_0/1counter_0/an2v0x3_3/zn 3seg_0/2seg_0/1counter_0/an2v0x3_3/b 2.4fF
C565 gnd 3seg_0/2seg_0/1counter_0/tf_0/xor2v0x05_0/a 8.1fF
C566 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_2/a 34.4fF
C567 decoder_0/or2v0x3_0/zn decoder_0/or2v0x3_0/z 2.3fF
C568 3seg_0/2seg_0/or3v0x3_0/a 3seg_0/2seg_0/totdiff3_0/mux_0/a0 2.3fF
C569 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_4/z 9.2fF
C570 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_3/z 12.6fF
C571 gnd 3seg_0/firseg_0/decoder_0/d6 48.5fF
C572 3seg_0/firseg_0/comp_0/an2v0x2_3/z vdd 9.1fF
C573 vdd 3seg_0/firseg_0/comp_0/an3v0x2_2/zn 4.9fF
C574 gnd 3seg_0/firseg_0/3_bitmux_0/mxn2v0x1_0/w_n4_n4# 76.0fF
C575 vdd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/d 9.8fF
C576 3seg_0/2seg_0/1counter_0/bf1v0x4_2/a 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/ci 2.1fF
C577 decoder_0/d1 decoder_0/or2v0x3_3/z 2.2fF
C578 3seg_0/2seg_0/totdiff3_0/diff2_2/xnr2v8x05_0/bn vdd 14.4fF
C579 3seg_0/firseg_0/comp_0/or3v0x2_0/zn 3seg_0/firseg_0/decoder_0/b0 3.3fF
C580 3seg_0/firseg_0/3_bitmux_0/o0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/zn 4.3fF
C581 3seg_0/2seg_0/1counter_0/or2v0x3_0/z 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/d 3.1fF
C582 vdd 3seg_0/firseg_0/comp_0/an3v0x2_3/zn 10.7fF
C583 gnd 3seg_0/2seg_0/an2v0x3_0/z 19.2fF
C584 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_1/zn 8.9fF
C585 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_8/zn 9.0fF
C586 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/an 6.8fF
C587 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_1/zn vdd 8.8fF
C588 decoder_0/d2 decoder_0/or2v0x3_0/z 2.2fF
C589 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/cn 3seg_0/2seg_0/totdiff3_0/mux_0/a2 4.1fF
C590 3seg_0/firseg_0/decoder_0/d0 gnd 7.6fF
C591 vdd decoder_0/or2v0x3_3/zn 12.7fF
C592 vdd 3seg_0/2seg_0/totdiff3_0/diff2_2/xor2v2x2_0/bn 17.7fF
C593 3seg_0/firseg_0/comp_0/an2v0x2_3/zn gnd 8.9fF
C594 3seg_0/2seg_0/1counter_0/an2v0x3_3/zn vdd 13.3fF
C595 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/cn 2.3fF
C596 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xnr2v8x05_0/zn 15.0fF
C597 gnd 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_2/a 25.9fF
C598 3seg_0/2seg_0/totdiff3_0/mux_0/b0 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an 3.9fF
C599 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/a 61.1fF
C600 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/or2v0x3_0/zn 9.0fF
C601 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_2/zn 8.9fF
C602 vdd 3seg_0/firseg_0/decoder_0/d5 21.8fF
C603 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/bn 11.2fF
C604 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/a2 36.6fF
C605 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/iz 3seg_0/2seg_0/totdiff3_0/diff2_2/xor3v1x2_0/bn 2.4fF
C606 3seg_0/2seg_0/totdiff3_0/mux_0/b1 3seg_0/2seg_0/totdiff3_0/mux_0/a1 39.4fF
C607 gnd 3seg_0/firseg_0/comp_0/an3v0x2_3/z 10.6fF
C608 3seg_0/2seg_0/ud 3seg_0/2seg_0/totdiff3_0/mux_0/mxn2v0x1_0/w_n4_n4# 30.3fF
C609 gnd 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/an 9.2fF
C610 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_1/a 31.8fF
C611 3seg_0/2seg_0/1counter_0/tf_1/dfnt1v0x2_0/n4 vdd 8.9fF
C612 vdd decoder_0/b2 16.7fF
C613 decoder_0/d1 decoder_0/or2v0x3_3/zn 3.7fF
C614 vdd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor3v1x2_0/iz 15.8fF
C615 3seg_0/2seg_0/1counter_0/or2v0x3_0/z vdd 11.4fF
C616 vdd 3seg_0/firseg_0/decoder_0/or2v0x3_3/zn 12.7fF
C617 vdd 3seg_0/2seg_0/or3v0x3_0/c 10.0fF
C618 gnd 3seg_0/firseg_0/decoder_0/or2v0x3_0/z 10.3fF
C619 gnd 3seg_0/2seg_0/an2v0x3_0/zn 9.5fF
C620 gnd 3seg_0/2seg_0/1counter_0/an2v0x3_2/z 16.1fF
C621 3seg_0/2seg_0/totdiff3_0/mux_0/a1 3seg_0/2seg_0/totdiff3_0/diff2_1/xor3v1x2_0/cn 4.1fF
C622 3seg_0/2seg_0/1counter_0/or2v0x3_1/z vdd 11.7fF
C623 gnd 3seg_0/firseg_0/3_bitmux_0/o0 60.8fF
C624 3seg_0/firseg_0/decoder_0/or2v0x3_3/z 3seg_0/firseg_0/decoder_0/d1 2.2fF
C625 gnd 3seg_0/2seg_0/totdiff3_0/diff2_1/xor2v2x2_0/an 21.6fF
C626 gnd 3seg_0/2seg_0/totdiff3_0/diff2_0/xor2v2x2_0/an 21.6fF
C627 vdd 3seg_0/2seg_0/totdiff3_0/mux_0/b2 3.1fF
C628 vdd 3seg_0/2seg_0/1counter_0/tf_0/dfnt1v0x2_0/n2 12.4fF
C629 decoder_0/or2v0x3_4/zn decoder_0/d6 2.1fF
C630 gnd 3seg_0/firseg_0/comp_0/an3v0x2_2/z 10.7fF
C631 3seg_0/firseg_0/comp_0/an3v0x2_2/w_n4_32# 3seg_0/firseg_0/comp_0/an3v0x2_1/a 8.3fF
C632 3seg_0/2seg_0/1counter_0/tf_2/dfnt1v0x2_0/d 3seg_0/2seg_0/1counter_0/tf_2/xor2v0x05_0/bn 2.8fF
C633 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z gnd 39.5fF
C634 decoder_0/d2 gnd! 12.7fF
C635 decoder_0/d0 gnd! 5.5fF
C636 decoder_0/d4 gnd! 25.7fF
C637 decoder_0/b0 gnd! 75.5fF
C638 vdd gnd! 910.6fF
C639 decoder_0/d5 gnd! 18.7fF
C640 decoder_0/d1 gnd! 15.2fF
C641 decoder_0/b1 gnd! 43.0fF
C642 decoder_0/d6 gnd! 2.7fF
C643 gnd gnd! 683.7fF
C644 decoder_0/d3 gnd! 17.6fF
C645 3seg_0/firseg_0/decoder_0/d2 gnd! 12.7fF
C646 3seg_0/firseg_0/decoder_0/d0 gnd! 5.5fF
C647 3seg_0/firseg_0/decoder_0/d4 gnd! 25.7fF
C648 3seg_0/firseg_0/decoder_0/d5 gnd! 18.7fF
C649 3seg_0/firseg_0/decoder_0/d1 gnd! 15.2fF
C650 3seg_0/firseg_0/decoder_0/d6 gnd! 2.7fF
C651 3seg_0/firseg_0/decoder_0/d3 gnd! 17.6fF
C652 decoder_0/b2 gnd! 45.2fF
C653 3seg_0/firseg_0/decoder_0/b0 gnd! 45.1fF
C654 3seg_0/firseg_0/comp_0/nr3v0x2_0/a gnd! 8.6fF
C655 3seg_0/firseg_0/3_bitmux_0/o0 gnd! 118.1fF
C656 3seg_0/firseg_0/out gnd! 43.1fF
C657 3seg_0/firseg_0/3_bitmux_0/o1 gnd! 73.8fF
C658 3seg_0/firseg_0/decoder_0/b1 gnd! 20.6fF
C659 3seg_0/firseg_0/3_bitmux_0/o2 gnd! 28.4fF
C660 3seg_0/firseg_0/decoder_0/b2 gnd! 36.6fF
C661 3seg_0/2seg_0/1counter_0/bf1v0x4_0/z gnd! 58.3fF
C662 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/b gnd! 2.9fF
C663 3seg_0/2seg_0/totdiff3_0/diff2_1/in_c gnd! 37.1fF
C664 3seg_0/2seg_0/totdiff3_0/diff2_0/an2v0x2_0/z gnd! 5.0fF
C665 3seg_0/2seg_0/1counter_0/bf1v0x4_1/z gnd! 39.5fF
C666 3seg_0/2seg_0/totdiff3_0/mux_0/a1 gnd! 28.9fF
C667 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/b gnd! 2.9fF
C668 3seg_0/2seg_0/totdiff3_0/diff2_2/in_c gnd! 36.8fF
C669 3seg_0/2seg_0/totdiff3_0/diff2_1/an2v0x2_0/z gnd! 5.0fF
C670 3seg_0/2seg_0/totdiff3_0/diff2_1/in_2c gnd! 29.6fF
C671 3seg_0/2seg_0/1counter_0/bf1v0x4_2/z gnd! 36.9fF
C672 3seg_0/2seg_0/totdiff3_0/mux_0/a2 gnd! 38.7fF
C673 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/b gnd! 2.9fF
C674 3seg_0/2seg_0/totdiff3_0/diff2_2/an2v0x2_0/z gnd! 5.0fF
C675 3seg_0/2seg_0/totdiff3_0/diff2_2/in_2c gnd! 34.8fF
C676 3seg_0/2seg_0/or3v0x3_0/a gnd! 68.8fF
C677 3seg_0/2seg_0/totdiff3_0/mux_0/b0 gnd! 47.5fF
C678 3seg_0/2seg_0/ud gnd! 52.0fF
C679 3seg_0/2seg_0/totdiff3_0/mux_0/a0 gnd! 99.1fF
C680 3seg_0/2seg_0/or3v0x3_0/b gnd! 71.7fF
C681 3seg_0/2seg_0/totdiff3_0/mux_0/b1 gnd! 87.1fF
C682 3seg_0/2seg_0/or3v0x3_0/c gnd! 52.7fF
C683 3seg_0/2seg_0/totdiff3_0/mux_0/b2 gnd! 24.6fF
C684 3seg_0/2seg_0/iv1v0x3_0/z gnd! 6.0fF
C685 3seg_0/2seg_0/1counter_0/or2v0x3_1/a gnd! 2.9fF
C686 3seg_0/2seg_0/1counter_0/an2v0x3_3/b gnd! 17.2fF
C687 3seg_0/2seg_0/1counter_0/bf1v0x4_2/a gnd! 2.3fF
C688 3seg_0/2seg_0/1counter_0/an2v0x3_2/z gnd! 4.6fF
C689 3seg_0/2seg_0/1counter_0/bf1v0x4_1/a gnd! 6.2fF
C690 3seg_0/2seg_0/1counter_0/an2v0x3_2/b gnd! 21.1fF
C691 3seg_0/2seg_0/1counter_0/an2v0x3_1/a gnd! 5.9fF
