* Spice description of mx3_x2
* Spice driver version 134999461
* Date 21/07/2007 at 19:29:40
* sxlib 0.13um values
.subckt mx3_x2 cmd0 cmd1 i0 i1 i2 q vdd vss
Mtr_00001 vss   cmd1  sig5  vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00002 sig12 cmd0  vss   vss n  L=0.12U  W=0.32U  AS=0.0848P   AD=0.0848P   PS=1.17U   PD=1.17U
Mtr_00003 sig2  i1    sig3  vss n  L=0.12U  W=0.65U  AS=0.17225P  AD=0.17225P  PS=1.83U   PD=1.83U
Mtr_00004 sig3  cmd1  sig4  vss n  L=0.12U  W=0.65U  AS=0.17225P  AD=0.17225P  PS=1.83U   PD=1.83U
Mtr_00005 sig4  sig5  sig1  vss n  L=0.12U  W=0.65U  AS=0.17225P  AD=0.17225P  PS=1.83U   PD=1.83U
Mtr_00006 sig1  i2    sig2  vss n  L=0.12U  W=0.65U  AS=0.17225P  AD=0.17225P  PS=1.83U   PD=1.83U
Mtr_00007 vss   cmd0  sig2  vss n  L=0.12U  W=0.65U  AS=0.17225P  AD=0.17225P  PS=1.83U   PD=1.83U
Mtr_00008 sig11 sig12 vss   vss n  L=0.12U  W=0.65U  AS=0.17225P  AD=0.17225P  PS=1.83U   PD=1.83U
Mtr_00009 sig4  i0    sig11 vss n  L=0.12U  W=0.65U  AS=0.17225P  AD=0.17225P  PS=1.83U   PD=1.83U
Mtr_00010 vss   sig4  q     vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00011 sig18 sig5  sig4  vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00012 vdd   sig12 sig17 vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00013 sig19 cmd0  vdd   vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00014 sig4  i0    sig19 vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00015 sig17 i1    sig18 vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00016 sig16 i2    sig17 vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00017 sig4  cmd1  sig16 vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00018 q     sig4  vdd   vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00019 sig5  cmd1  vdd   vdd p  L=0.12U  W=0.76U  AS=0.2014P   AD=0.2014P   PS=2.05U   PD=2.05U
Mtr_00020 vdd   cmd0  sig12 vdd p  L=0.12U  W=0.76U  AS=0.2014P   AD=0.2014P   PS=2.05U   PD=2.05U
C14 cmd0  vss   0.823f
C9  cmd1  vss   0.887f
C15 i0    vss   0.713f
C8  i1    vss   0.393f
C10 i2    vss   0.338f
C13 q     vss   0.980f
C12 sig12 vss   0.821f
C17 sig17 vss   0.344f
C2  sig2  vss   0.344f
C4  sig4  vss   1.569f
C5  sig5  vss   0.787f
.ends
