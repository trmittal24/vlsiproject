* Spice description of nd3_x05
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:10
*
.subckt nd3_x05 a b c vdd vss z 
M1  z     c     vdd   vdd p  L=0.13U  W=0.605U AS=0.160325P AD=0.160325P PS=1.74U   PD=1.74U  
M3  z     a     vdd   vdd p  L=0.13U  W=0.605U AS=0.160325P AD=0.160325P PS=1.74U   PD=1.74U  
M2  vdd   b     z     vdd p  L=0.13U  W=0.605U AS=0.160325P AD=0.160325P PS=1.74U   PD=1.74U  
M4  n2    c     z     vss n  L=0.13U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U  
M5  n1    b     n2    vss n  L=0.13U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U  
M6  vss   a     n1    vss n  L=0.13U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U  
C8  vdd   vss   1.476f
C7  a     vss   0.726f
C6  c     vss   1.097f
C5  b     vss   0.757f
C2  z     vss   2.282f
.ends
