* Spice description of nao2o22_x4
* Spice driver version 134999461
* Date 31/05/2007 at 10:38:17
* ssxlib 0.13um values
.subckt nao2o22_x4 i0 i1 i2 i3 nq vdd vss
Mtr_00001 sig9  sig1  vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00002 nq    sig9  vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00003 vss   sig9  nq    vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00004 sig2  i3    vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00005 vss   i2    sig2  vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00006 sig2  i0    sig1  vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00007 sig1  i1    sig2  vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00008 vdd   sig1  sig9  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00009 vdd   sig9  nq    vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
Mtr_00010 nq    sig9  vdd   vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
Mtr_00011 sig11 i0    vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00012 sig12 i3    sig1  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00013 vdd   i2    sig12 vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00014 sig1  i1    sig11 vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
C4  i0    vss   0.660f
C5  i1    vss   0.688f
C7  i2    vss   0.660f
C6  i3    vss   0.688f
C8  nq    vss   0.771f
C1  sig1  vss   1.098f
C2  sig2  vss   0.345f
C9  sig9  vss   0.702f
.ends
