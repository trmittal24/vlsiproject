* Sat Aug 27 19:34:31 CEST 2005
.subckt nd2v4x4 a b vdd vss z 
*SPICE circuit <nd2v4x4> from XCircuit v3.20

m1 n1 a vss vss n w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m2 z a vdd vdd p w=62u l=2u ad='62u*5u+12p' as='62u*5u+12p' pd='62u*2+14u' ps='62u*2+14u'
m3 z b n1 vss n w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m4 z b vdd vdd p w=62u l=2u ad='62u*5u+12p' as='62u*5u+12p' pd='62u*2+14u' ps='62u*2+14u'
.ends
