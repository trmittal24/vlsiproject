* Tue Aug 10 11:21:07 CEST 2004
.subckt bf1_w05 a vdd vss z 
*SPICE circuit <bf1_w05> from XCircuit v3.10

m1 an a vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m2 an a vdd vdd p w=9u l=2u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m3 z an vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m4 z an vdd vdd p w=9u l=2u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
.ends
