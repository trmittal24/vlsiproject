* Spice description of oai21v0x05
* Spice driver version 134999461
* Date 17/05/2007 at  9:30:05
* vsclib 0.13um values
.subckt oai21v0x05 a1 a2 b vdd vss z
M01 vdd   a1    n2    vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M02 sig1  a1    vss   vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M03 n2    a2    z     vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M04 vss   a2    sig1  vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M05 z     b     vdd   vdd p  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M06 sig1  b     z     vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
C6  a1    vss   0.357f
C4  a2    vss   0.461f
C5  b     vss   0.466f
C1  sig1  vss   0.226f
C2  z     vss   0.818f
.ends
