* Mon Aug 16 14:10:59 CEST 2004
.subckt nd2v0x05 a b vdd vss z 
*SPICE circuit <nd2v0x05> from XCircuit v3.10

m1 n1 a vss vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m2 z a vdd vdd p w=8u l=2u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
m3 z b n1 vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m4 z b vdd vdd p w=8u l=2u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
.ends
