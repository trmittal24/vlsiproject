magic
tech scmos
timestamp 1523003210
<< nwell >>
rect -282 75 -268 85
<< metal1 >>
rect -221 150 114 157
rect -277 131 -259 135
rect -277 102 -273 131
rect 7 115 62 118
rect -275 85 -215 90
rect -282 78 -215 85
rect -371 75 -215 78
rect 46 77 107 91
rect -371 69 -280 75
rect -273 73 -215 75
rect -76 69 134 77
rect 138 69 153 77
rect -292 55 -284 56
rect 5 55 14 56
rect -288 51 -284 55
rect 7 51 14 55
rect -478 46 -467 47
rect -478 43 -477 46
rect -473 43 -467 46
rect -403 44 -402 46
rect -407 36 -402 44
rect -177 42 -175 46
rect 116 46 121 47
rect -111 38 -107 44
rect 118 43 121 46
rect -111 35 -108 38
rect -268 23 -264 30
rect -15 22 -12 28
rect 28 22 32 28
rect -373 5 -282 14
rect -84 11 145 13
rect -271 -6 -211 11
rect -84 5 150 11
rect 50 -11 150 5
rect -268 -25 -264 -20
rect -268 -29 -256 -25
rect 29 -28 71 -25
rect 25 -29 71 -28
rect 129 -29 133 -24
rect 104 -68 123 -67
rect -220 -75 123 -68
<< metal2 >>
rect -9 123 99 126
rect -9 117 -6 123
rect -260 114 -59 117
rect -38 114 -6 117
rect -305 106 -224 109
rect -421 55 -352 59
rect -421 45 -417 55
rect -355 48 -352 55
rect -305 49 -302 106
rect -277 87 -273 98
rect -292 84 -273 87
rect -292 55 -288 84
rect -9 49 -6 114
rect 3 55 6 114
rect -473 42 -417 45
rect -403 44 -388 47
rect -355 45 -322 48
rect -392 39 -388 44
rect -326 39 -322 45
rect -198 42 -181 46
rect -177 42 -131 45
rect -107 44 -59 47
rect -198 39 -195 42
rect -392 37 -355 39
rect -392 35 -359 37
rect -326 36 -195 39
rect -134 38 -131 42
rect -63 40 -59 44
rect -134 35 -67 38
rect 101 42 114 45
rect -134 34 -131 35
rect -70 29 -67 35
rect 101 29 104 42
rect -70 26 104 29
rect -311 -31 -308 24
rect -268 -16 -265 19
rect -311 -34 -219 -31
rect -15 -32 -12 18
rect 25 -24 28 22
rect -15 -35 102 -32
rect -259 -57 -256 -46
rect 41 -57 44 -35
rect -259 -60 -3 -57
rect 18 -60 44 -57
rect 62 -62 65 -46
rect 140 -62 144 -53
rect 62 -65 144 -62
<< m2contact >>
rect 99 123 103 127
rect -264 114 -260 118
rect 3 114 7 118
rect -224 105 -220 109
rect -277 98 -273 102
rect -292 51 -288 55
rect 3 51 7 55
rect -477 42 -473 46
rect -407 44 -403 48
rect -305 45 -301 49
rect -181 42 -177 46
rect -111 44 -107 48
rect -9 45 -5 49
rect 114 42 118 46
rect -359 33 -355 37
rect -63 36 -59 40
rect -312 24 -308 28
rect -268 19 -264 23
rect -16 18 -12 22
rect 28 18 32 22
rect -268 -20 -264 -16
rect 25 -28 29 -24
rect -219 -34 -215 -30
rect 102 -35 106 -31
rect -260 -46 -256 -42
rect 61 -46 65 -42
rect 140 -53 144 -49
use ../pharosc_8.4/magic/cells/vsclib/an2v0x3  an2v0x3_3
timestamp 1522990558
transform -1 0 -217 0 -1 157
box -4 -4 60 76
use ../pharosc_8.4/magic/cells/vsclib/an2v0x3  an2v0x3_0
timestamp 1522990558
transform -1 0 105 0 -1 157
box -4 -4 60 76
use tf  tf_2
timestamp 1522990558
transform 1 0 -589 0 1 1
box 0 0 224 80
use ../pharosc_8.4/magic/cells/vsclib/or2v0x3  or2v0x3_1
timestamp 1522990558
transform 1 0 -361 0 1 5
box -4 -4 68 76
use tf  tf_1
timestamp 1522990558
transform 1 0 -293 0 1 1
box 0 0 224 80
use ../pharosc_8.4/magic/cells/vsclib/or2v0x3  or2v0x3_0
timestamp 1522990558
transform 1 0 -65 0 1 5
box -4 -4 68 76
use tf  tf_0
timestamp 1522990558
transform 1 0 3 0 1 1
box 0 0 224 80
use ../pharosc_8.4/magic/cells/vsclib/an2v0x3  an2v0x3_2
timestamp 1522990558
transform -1 0 -213 0 -1 -3
box -4 -4 60 76
use ../pharosc_8.4/magic/cells/vsclib/an2v0x3  an2v0x3_1
timestamp 1522990558
transform -1 0 108 0 -1 -3
box -4 -4 60 76
use ../pharosc_8.4/magic/cells/vsclib/iv1v0x3  iv1v0x3_0
timestamp 1522990558
transform -1 0 148 0 -1 -3
box -4 -4 36 76
<< end >>
