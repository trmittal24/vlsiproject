* Mon Aug 16 14:10:59 CEST 2004
.subckt nd2v0x4 a b vdd vss z 
*SPICE circuit <nd2v0x4> from XCircuit v3.10

m1 n1 a vss vss n w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m2 z a vdd vdd p w=48u l=2.3636u ad='48u*5u+12p' as='48u*5u+12p' pd='48u*2+14u' ps='48u*2+14u'
m3 z b n1 vss n w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m4 z b vdd vdd p w=48u l=2.3636u ad='48u*5u+12p' as='48u*5u+12p' pd='48u*2+14u' ps='48u*2+14u'
.ends
