* Fri Apr  8 11:37:06 CEST 2005
.subckt aoi22v0x4 a1 a2 b1 b2 vdd vss z 
*SPICE circuit <aoi22v0x4> from XCircuit v3.20

m1 n1 b1 vss vss n w=50u l=2u ad='50u*5u+12p' as='50u*5u+12p' pd='50u*2+14u' ps='50u*2+14u'
m2 z b1 n3 vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
m3 n3 a1 vdd vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
m4 n3 a2 vdd vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
m5 n2 a1 vss vss n w=50u l=2u ad='50u*5u+12p' as='50u*5u+12p' pd='50u*2+14u' ps='50u*2+14u'
m6 z b2 n1 vss n w=50u l=2u ad='50u*5u+12p' as='50u*5u+12p' pd='50u*2+14u' ps='50u*2+14u'
m7 z a2 n2 vss n w=50u l=2u ad='50u*5u+12p' as='50u*5u+12p' pd='50u*2+14u' ps='50u*2+14u'
m8 z b2 n3 vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
.ends
