* Wed Apr  5 08:55:15 CEST 2006
.subckt bf1v2x1 a vdd vss z 
*SPICE circuit <bf1v2x1> from XCircuit v3.20

m1 an a vss vss n w=7u l=2.3636u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m2 an a vdd vdd p w=14u l=2.3636u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m3 z an vss vss n w=9u l=2.3636u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m4 z an vdd vdd p w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
.ends
