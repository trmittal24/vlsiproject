* Tue Feb 27 17:14:04 CET 2007
.subckt nd3v5x4 a b c vdd vss z
*SPICE circuit <nd3v5x4> from XCircuit v3.4 rev 26

m1 z c vdd vdd p w=60u l=2u ad='60u*5u+12p' as='60u*5u+12p' pd='60u*2+14u' ps='60u*2+14u'
m2 z a vdd vdd p w=60u l=2u ad='60u*5u+12p' as='60u*5u+12p' pd='60u*2+14u' ps='60u*2+14u'
m3 n1 a vss vss n w=60u l=2u ad='60u*5u+12p' as='60u*5u+12p' pd='60u*2+14u' ps='60u*2+14u'
m4 n2 b n1 vss n w=60u l=2u ad='60u*5u+12p' as='60u*5u+12p' pd='60u*2+14u' ps='60u*2+14u'
m5 z c n2 vss n w=60u l=2u ad='60u*5u+12p' as='60u*5u+12p' pd='60u*2+14u' ps='60u*2+14u'
m6 z b vdd vdd p w=60u l=2u ad='60u*5u+12p' as='60u*5u+12p' pd='60u*2+14u' ps='60u*2+14u'
.ends
