* Mon Aug 16 14:10:56 CEST 2004
.subckt an4v0x1 a b c d vdd vss z 
*SPICE circuit <an4v0x1> from XCircuit v3.10

m1 zn a vdd vdd p w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m2 zn b vdd vdd p w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m3 zn c vdd vdd p w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m4 zn d n3 vss n w=16u l=2.3636u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m5 n3 c n2 vss n w=16u l=2.3636u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m6 n2 b n1 vss n w=16u l=2.3636u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m7 z zn vss vss n w=9u l=2.3636u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m8 z zn vdd vdd p w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m9 zn d vdd vdd p w=13u l=2.3636u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m10 n1 a vss vss n w=16u l=2.3636u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
.ends
