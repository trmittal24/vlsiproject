* Spice description of tie_x0
* Spice driver version 134999461
* Date 31/05/2007 at 10:40:36
* ssxlib 0.13um values
.subckt tie_x0 vdd vss
.ends
