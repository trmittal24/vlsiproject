* Tue Feb 20 08:57:11 CET 2007
.subckt aoi21v0x1 a1 a2 b vdd vss z
*SPICE circuit <aoi21v0x1> from XCircuit v3.4 rev 26

m1 n1 a2 vdd vdd p w=26u l=2.3636u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m2 n1 a1 vdd vdd p w=26u l=2.3636u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m3 n2 a1 vss vss n w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m4 z b vss vss n w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m5 z a2 n2 vss n w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m6 z b n1 vdd p w=26u l=2.3636u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
.ends
