* Sat Aug 27 22:10:03 CEST 2005
.subckt iv1v4x3 a vdd vss z 
*SPICE circuit <iv1v4x3> from XCircuit v3.20

m1 z a vss vss n w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m2 z a vdd vdd p w=48u l=2.3636u ad='48u*5u+12p' as='48u*5u+12p' pd='48u*2+14u' ps='48u*2+14u'
.ends
