magic
tech scmos
timestamp 1521974529
use xor3v1x2  xor3v1x2_0
timestamp 1521974529
transform 1 0 4 0 1 4
box -4 -4 172 76
<< end >>
