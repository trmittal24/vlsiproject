* Tue Dec 14 18:00:58 CET 2004
.subckt xooi21v0x2 a1 a2 b vdd vss z 
*SPICE circuit <xooi21v0x2> from XCircuit v3.20

m1 an a1 vss vss n w=24u l=2u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m2 an a2 vss vss n w=24u l=2u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m3 n1 a1 vdd vdd p w=72u l=2u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
m4 an a2 n1 vdd p w=72u l=2u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
m5 n2 bn vdd vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m6 z b an vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m7 bn b vss vss n w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m8 z an bn vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m9 bn b vdd vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m10 z bn an vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m11 z an n2 vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
.ends
