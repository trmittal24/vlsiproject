* Fri Mar 31 22:05:19 CEST 2006
.subckt an2v2x2 a b vdd vss z 
*SPICE circuit <an2v2x2> from XCircuit v3.20

m1 z zn vdd vdd p w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m2 z zn vss vss n w=14u l=2u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m3 n1 a vss vss n w=14u l=2u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m4 zn a vdd vdd p w=17u l=2u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m5 zn b n1 vss n w=14u l=2u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m6 zn b vdd vdd p w=17u l=2u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
.ends
