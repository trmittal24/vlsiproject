* Spice description of bf1v2x3
* Spice driver version 134999461
* Date 17/05/2007 at  9:05:32
* wsclib 0.13um values
.subckt bf1v2x3 a vdd vss z
M01 05    a     vdd   vdd p  L=0.12U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U
M02 05    a     vss   vss n  L=0.12U  W=0.605U AS=0.160325P AD=0.160325P PS=1.74U   PD=1.74U
M03 z     05    vdd   vdd p  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
M04 vdd   05    z     vdd p  L=0.12U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U
M05 vss   05    z     vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
C3  05    vss   0.541f
C4  a     vss   0.472f
C2  z     vss   0.637f
.ends
