* Sun Nov 28 12:41:02 CET 2004
.subckt nr2av1x05 a b vdd vss z 
*SPICE circuit <nr2av1x05> from XCircuit v3.20

m1 an a vss vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m2 an a vdd vdd p w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m3 z an vss vss n w=8u l=2.3636u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
m4 n1 an vdd vdd p w=15u l=2.3636u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m5 z b vss vss n w=8u l=2.3636u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
m6 z b n1 vdd p w=15u l=2.3636u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
.ends
