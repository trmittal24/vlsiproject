* Mon Aug 16 14:10:59 CEST 2004
.subckt nd4v0x3 a b c d vdd vss z 
*SPICE circuit <nd4v0x3> from XCircuit v3.10

m1 z a vdd vdd p w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m2 z b vdd vdd p w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m3 z c vdd vdd p w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m4 z d vdd vdd p w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m5 n1 a vss vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m6 n2 b n1 vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m7 n3 c n2 vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m8 z d n3 vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
.ends
