* Mon Apr 16 10:17:40 CEST 2007
.subckt xnr2v0x4 a b vdd vss z
*SPICE circuit <xnr2v0x4> from XCircuit v3.4 rev 26

m1 n1 bn vdd vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
m2 z b an vdd p w=75u l=2u ad='75u*5u+12p' as='75u*5u+12p' pd='75u*2+14u' ps='75u*2+14u'
m3 bn b vss vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m4 an a vss vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m5 z an bn vss n w=38u l=2u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m6 an a vdd vdd p w=75u l=2u ad='75u*5u+12p' as='75u*5u+12p' pd='75u*2+14u' ps='75u*2+14u'
m7 bn b vdd vdd p w=75u l=2u ad='75u*5u+12p' as='75u*5u+12p' pd='75u*2+14u' ps='75u*2+14u'
m8 z bn an vss n w=36u l=2u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
m9 z an n1 vdd p w=112u l=2u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
.ends
