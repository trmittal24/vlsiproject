* SPICE3 file created from comp.ext - technology: scmos

.include t14y_tsmc_025_level3.txt

.option scale=1u

M1000 nr2v0x2_0_a_11_39# nr2v0x2_0_a iv1v0x4_2_vdd iv1v0x4_2_vdd pfet w=27 l=2
+ ad=135 pd=64 as=3890 ps=1322 
M1001 nr2v0x2_0_z an2v0x2_1_z nr2v0x2_0_a_11_39# iv1v0x4_2_vdd pfet w=27 l=2
+ ad=216 pd=70 as=0 ps=0 
M1002 nr2v0x2_0_a_28_39# an2v0x2_1_z nr2v0x2_0_z iv1v0x4_2_vdd pfet w=27 l=2
+ ad=135 pd=64 as=0 ps=0 
M1003 iv1v0x4_2_vdd nr2v0x2_0_a nr2v0x2_0_a_28_39# iv1v0x4_2_vdd pfet w=27 l=2
+ ad=0 pd=0 as=0 ps=0 
M1004 nr2v0x2_0_z nr2v0x2_0_a iv1v0x4_0_vss iv1v0x4_0_vss nfet w=15 l=2
+ ad=120 pd=46 as=2273 ps=830 
M1005 iv1v0x4_0_vss an2v0x2_1_z nr2v0x2_0_z iv1v0x4_0_vss nfet w=15 l=2
+ ad=0 pd=0 as=0 ps=0 
M1006 iv1v0x4_2_vdd or3v0x2_1_zn or3v0x2_1_z iv1v0x4_2_vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1007 or3v0x2_1_a_24_38# iv1v0x4_2_z iv1v0x4_2_vdd iv1v0x4_2_vdd pfet w=22 l=2
+ ad=110 pd=54 as=0 ps=0 
M1008 or3v0x2_1_a_31_38# or3v0x2_0_c or3v0x2_1_a_24_38# iv1v0x4_2_vdd pfet w=22 l=2
+ ad=110 pd=54 as=0 ps=0 
M1009 or3v0x2_1_zn or3v0x2_1_c or3v0x2_1_a_31_38# iv1v0x4_2_vdd pfet w=22 l=2
+ ad=167 pd=60 as=0 ps=0 
M1010 or3v0x2_1_a_48_38# or3v0x2_1_c or3v0x2_1_zn iv1v0x4_2_vdd pfet w=19 l=2
+ ad=95 pd=48 as=0 ps=0 
M1011 or3v0x2_1_a_55_38# or3v0x2_0_c or3v0x2_1_a_48_38# iv1v0x4_2_vdd pfet w=19 l=2
+ ad=95 pd=48 as=0 ps=0 
M1012 iv1v0x4_2_vdd iv1v0x4_2_z or3v0x2_1_a_55_38# iv1v0x4_2_vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1013 iv1v0x4_0_vss or3v0x2_1_zn or3v0x2_1_z iv1v0x4_0_vss nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1014 or3v0x2_1_zn iv1v0x4_2_z iv1v0x4_0_vss iv1v0x4_0_vss nfet w=8 l=2
+ ad=116 pd=62 as=0 ps=0 
M1015 iv1v0x4_0_vss or3v0x2_0_c or3v0x2_1_zn iv1v0x4_0_vss nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1016 or3v0x2_1_zn or3v0x2_1_c iv1v0x4_0_vss iv1v0x4_0_vss nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1017 iv1v0x4_2_vdd an2v0x2_1_zn an2v0x2_1_z iv1v0x4_2_vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1018 an2v0x2_1_zn an2v0x2_0_z iv1v0x4_2_vdd iv1v0x4_2_vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1019 iv1v0x4_2_vdd an2v0x2_1_b an2v0x2_1_zn iv1v0x4_2_vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1020 iv1v0x4_0_vss an2v0x2_1_zn an2v0x2_1_z iv1v0x4_0_vss nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1021 an2v0x2_1_a_24_13# an2v0x2_0_z iv1v0x4_0_vss iv1v0x4_0_vss nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1022 an2v0x2_1_zn an2v0x2_1_b an2v0x2_1_a_24_13# iv1v0x4_0_vss nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1023 iv1v0x4_2_vdd an2v0x2_0_zn an2v0x2_0_z iv1v0x4_2_vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1024 an2v0x2_0_zn an2v0x2_0_a iv1v0x4_2_vdd iv1v0x4_2_vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1025 iv1v0x4_2_vdd iv1v0x4_2_z an2v0x2_0_zn iv1v0x4_2_vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1026 iv1v0x4_0_vss an2v0x2_0_zn an2v0x2_0_z iv1v0x4_0_vss nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1027 an2v0x2_0_a_24_13# an2v0x2_0_a iv1v0x4_0_vss iv1v0x4_0_vss nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1028 an2v0x2_0_zn iv1v0x4_2_z an2v0x2_0_a_24_13# iv1v0x4_0_vss nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1029 iv1v0x4_2_z iv1v0x4_2_a iv1v0x4_2_vdd iv1v0x4_2_vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1030 iv1v0x4_2_vdd iv1v0x4_2_a iv1v0x4_2_z iv1v0x4_2_vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1031 iv1v0x4_2_z iv1v0x4_2_a iv1v0x4_0_vss iv1v0x4_0_vss nfet w=17 l=2
+ ad=118 pd=50 as=0 ps=0 
M1032 iv1v0x4_0_vss iv1v0x4_2_a iv1v0x4_2_z iv1v0x4_0_vss nfet w=11 l=2
+ ad=0 pd=0 as=0 ps=0 
M1033 iv1v0x4_2_vdd an2v0x2_3_zn nr2v0x2_0_a iv1v0x4_2_vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1034 an2v0x2_3_zn an2v0x2_2_z iv1v0x4_2_vdd iv1v0x4_2_vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1035 iv1v0x4_2_vdd or3v0x2_1_z an2v0x2_3_zn iv1v0x4_2_vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1036 iv1v0x4_0_vss an2v0x2_3_zn nr2v0x2_0_a iv1v0x4_0_vss nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1037 an2v0x2_3_a_24_13# an2v0x2_2_z iv1v0x4_0_vss iv1v0x4_0_vss nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1038 an2v0x2_3_zn or3v0x2_1_z an2v0x2_3_a_24_13# iv1v0x4_0_vss nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1039 iv1v0x4_2_vdd an2v0x2_2_zn an2v0x2_2_z iv1v0x4_2_vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1040 an2v0x2_2_zn an2v0x2_2_a iv1v0x4_2_vdd iv1v0x4_2_vdd pfet w=19 l=2
+ ad=152 pd=54 as=0 ps=0 
M1041 iv1v0x4_2_vdd or3v0x2_0_a an2v0x2_2_zn iv1v0x4_2_vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1042 iv1v0x4_0_vss an2v0x2_2_zn an2v0x2_2_z iv1v0x4_0_vss nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1043 an2v0x2_2_a_24_13# an2v0x2_2_a iv1v0x4_0_vss iv1v0x4_0_vss nfet w=13 l=2
+ ad=65 pd=36 as=0 ps=0 
M1044 an2v0x2_2_zn or3v0x2_0_a an2v0x2_2_a_24_13# iv1v0x4_0_vss nfet w=13 l=2
+ ad=77 pd=40 as=0 ps=0 
M1045 iv1v0x4_2_vdd or3v0x2_0_zn an2v0x2_1_b iv1v0x4_2_vdd pfet w=28 l=2
+ ad=0 pd=0 as=166 ps=70 
M1046 or3v0x2_0_a_24_38# or3v0x2_0_a iv1v0x4_2_vdd iv1v0x4_2_vdd pfet w=22 l=2
+ ad=110 pd=54 as=0 ps=0 
M1047 or3v0x2_0_a_31_38# or3v0x2_1_c or3v0x2_0_a_24_38# iv1v0x4_2_vdd pfet w=22 l=2
+ ad=110 pd=54 as=0 ps=0 
M1048 or3v0x2_0_zn or3v0x2_0_c or3v0x2_0_a_31_38# iv1v0x4_2_vdd pfet w=22 l=2
+ ad=167 pd=60 as=0 ps=0 
M1049 or3v0x2_0_a_48_38# or3v0x2_0_c or3v0x2_0_zn iv1v0x4_2_vdd pfet w=19 l=2
+ ad=95 pd=48 as=0 ps=0 
M1050 or3v0x2_0_a_55_38# or3v0x2_1_c or3v0x2_0_a_48_38# iv1v0x4_2_vdd pfet w=19 l=2
+ ad=95 pd=48 as=0 ps=0 
M1051 iv1v0x4_2_vdd or3v0x2_0_a or3v0x2_0_a_55_38# iv1v0x4_2_vdd pfet w=19 l=2
+ ad=0 pd=0 as=0 ps=0 
M1052 iv1v0x4_0_vss or3v0x2_0_zn an2v0x2_1_b iv1v0x4_0_vss nfet w=14 l=2
+ ad=0 pd=0 as=98 ps=42 
M1053 or3v0x2_0_zn or3v0x2_0_a iv1v0x4_0_vss iv1v0x4_0_vss nfet w=8 l=2
+ ad=116 pd=62 as=0 ps=0 
M1054 iv1v0x4_0_vss or3v0x2_1_c or3v0x2_0_zn iv1v0x4_0_vss nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1055 or3v0x2_0_zn or3v0x2_0_c iv1v0x4_0_vss iv1v0x4_0_vss nfet w=8 l=2
+ ad=0 pd=0 as=0 ps=0 
M1056 or3v0x2_0_c iv1v0x4_1_a iv1v0x4_2_vdd iv1v0x4_2_vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1057 iv1v0x4_2_vdd iv1v0x4_1_a or3v0x2_0_c iv1v0x4_2_vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1058 or3v0x2_0_c iv1v0x4_1_a iv1v0x4_0_vss iv1v0x4_0_vss nfet w=17 l=2
+ ad=118 pd=50 as=0 ps=0 
M1059 iv1v0x4_0_vss iv1v0x4_1_a or3v0x2_0_c iv1v0x4_0_vss nfet w=11 l=2
+ ad=0 pd=0 as=0 ps=0 
M1060 an2v0x2_0_a iv1v0x4_0_a iv1v0x4_2_vdd iv1v0x4_2_vdd pfet w=28 l=2
+ ad=224 pd=72 as=0 ps=0 
M1061 iv1v0x4_2_vdd iv1v0x4_0_a an2v0x2_0_a iv1v0x4_2_vdd pfet w=28 l=2
+ ad=0 pd=0 as=0 ps=0 
M1062 an2v0x2_0_a iv1v0x4_0_a iv1v0x4_0_vss iv1v0x4_0_vss nfet w=17 l=2
+ ad=118 pd=50 as=0 ps=0 
M1063 iv1v0x4_0_vss iv1v0x4_0_a an2v0x2_0_a iv1v0x4_0_vss nfet w=11 l=2
+ ad=0 pd=0 as=0 ps=0 
C0 or3v0x2_0_zn iv1v0x4_2_vdd 9.0fF
C1 iv1v0x4_2_vdd an2v0x2_2_zn 8.8fF
C2 iv1v0x4_1_a iv1v0x4_0_vss 8.9fF
C3 an2v0x2_0_zn iv1v0x4_2_vdd 8.8fF
C4 an2v0x2_0_z iv1v0x4_0_vss 9.8fF
C5 iv1v0x4_0_vss iv1v0x4_2_z 15.7fF
C6 iv1v0x4_2_vdd or3v0x2_1_z 13.7fF
C7 or3v0x2_1_zn iv1v0x4_0_vss 10.9fF
C8 iv1v0x4_2_a iv1v0x4_2_vdd 9.9fF
C9 or3v0x2_0_zn iv1v0x4_0_vss 10.9fF
C10 nr2v0x2_0_z iv1v0x4_2_vdd 4.3fF
C11 an2v0x2_2_zn iv1v0x4_0_vss 8.9fF
C12 an2v0x2_0_zn iv1v0x4_0_vss 8.9fF
C13 or3v0x2_1_c iv1v0x4_2_vdd 24.1fF
C14 an2v0x2_0_a iv1v0x4_2_vdd 13.4fF
C15 iv1v0x4_0_vss or3v0x2_1_z 15.0fF
C16 iv1v0x4_2_a iv1v0x4_0_vss 8.9fF
C17 nr2v0x2_0_z iv1v0x4_0_vss 5.5fF
C18 or3v0x2_0_c or3v0x2_0_zn 4.1fF
C19 an2v0x2_3_zn iv1v0x4_2_vdd 8.8fF
C20 or3v0x2_1_c iv1v0x4_0_vss 28.0fF
C21 an2v0x2_0_a iv1v0x4_0_vss 16.9fF
C22 an2v0x2_3_zn iv1v0x4_0_vss 8.9fF
C23 or3v0x2_0_c or3v0x2_1_c 2.9fF
C24 nr2v0x2_0_a iv1v0x4_2_vdd 9.1fF
C25 iv1v0x4_2_vdd or3v0x2_0_a 24.6fF
C26 nr2v0x2_0_a iv1v0x4_0_vss 20.8fF
C27 an2v0x2_2_z iv1v0x4_2_vdd 9.4fF
C28 iv1v0x4_0_a iv1v0x4_2_vdd 9.9fF
C29 or3v0x2_0_a iv1v0x4_0_vss 12.3fF
C30 iv1v0x4_2_vdd an2v0x2_2_a 6.6fF
C31 an2v0x2_1_b iv1v0x4_2_vdd 14.2fF
C32 an2v0x2_2_z iv1v0x4_0_vss 11.1fF
C33 iv1v0x4_0_a iv1v0x4_0_vss 8.9fF
C34 an2v0x2_2_a iv1v0x4_0_vss 5.5fF
C35 an2v0x2_1_b iv1v0x4_0_vss 5.9fF
C36 or3v0x2_0_c iv1v0x4_2_vdd 30.1fF
C37 an2v0x2_1_z iv1v0x4_2_vdd 22.0fF
C38 an2v0x2_1_zn iv1v0x4_2_vdd 8.8fF
C39 or3v0x2_0_c iv1v0x4_0_vss 34.3fF
C40 an2v0x2_1_z iv1v0x4_0_vss 8.7fF
C41 an2v0x2_1_zn iv1v0x4_0_vss 8.9fF
C42 iv1v0x4_2_vdd iv1v0x4_1_a 9.9fF
C43 an2v0x2_0_z iv1v0x4_2_vdd 10.7fF
C44 iv1v0x4_2_vdd iv1v0x4_2_z 37.6fF
C45 or3v0x2_1_zn iv1v0x4_2_vdd 9.0fF
C46 iv1v0x4_2_vdd 0 61.7fF

v_dd iv1v0x4_2_vdd 0 5
v_ss iv1v0x4_0_vss 0 0
v_gg_f iv1v0x4_1_a 0 PULSE(5 0 0 0.1n 0.1n 15n 30n)
v_gg_e iv1v0x4_2_a 0 PULSE(5 0 0 0.1n 0.1n 30n 60n)
v_gg_d iv1v0x4_0_a 0 PULSE(5 0 0 0.1n 0.1n 60n 120n)
v_gg_c or3v0x2_1_c 0 PULSE(5 0 0 0.1n 0.1n 120n 240n)
v_gg_b or3v0x2_0_a 0 PULSE(5 0 0 0.1n 0.1n 240n 480n)
v_gg_a an2v0x2_2_a 0 PULSE(5 0 0 0.1n 0.1n 480n 960n)

.control
 tran 0.01n 960n
 plot (an2v0x2_2_a + 5) (or3v0x2_0_a) (or3v0x2_1_c - 5) (iv1v0x4_0_a - 10) (iv1v0x4_2_a - 15) (iv1v0x4_1_a - 20) ( nr2v0x2_0_z - 25)
.endc

.end