* Spice description of vfeed4
* Spice driver version 134999461
* Date 22/07/2007 at 11:00:23
* vsxlib 0.13um values
.subckt vfeed4 vdd vss
.ends
