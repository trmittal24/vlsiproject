* Tue Feb 20 08:57:11 CET 2007
.subckt iv1v0x6 a vdd vss z
*SPICE circuit <iv1v0x6> from XCircuit v3.4 rev 26

m1 z a vss vss n w=54u l=2.3636u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m2 z a vdd vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
.ends
