* Spice description of vsstie
* Spice driver version 134999461
* Date 22/07/2007 at 11:00:32
* vsxlib 0.13um values
.subckt vsstie vdd vss z
M1  z     vdd   vdd   vdd p  L=0.12U  W=1.65U  AS=0.43725P  AD=0.43725P  PS=3.83U   PD=3.83U
M2  vss   vdd   z     vss n  L=0.12U  W=1.265U AS=0.335225P AD=0.335225P PS=3.06U   PD=3.06U
C1  z     vss   0.915f
.ends
