magic
tech scmos
timestamp 1523195521
<< polysilicon >>
rect 406 994 408 1008
<< metal1 >>
rect 11 1250 97 1255
rect 302 1176 327 1180
rect 70 1105 89 1112
rect 70 1001 77 1105
rect 323 1031 327 1176
rect 305 1027 327 1031
rect 407 1015 410 1218
rect 1032 1187 1035 1194
rect 406 1012 410 1015
rect 651 1184 1035 1187
rect 70 999 83 1001
rect 651 1000 654 1184
rect -21 994 83 999
rect -21 993 76 994
rect 629 982 650 986
rect 629 788 633 982
rect 1 766 77 775
rect 740 772 1010 773
rect 740 767 1034 772
rect 740 766 1010 767
rect 1025 685 1034 767
rect 905 586 1030 590
rect 1026 512 1030 586
rect 989 22 995 84
rect 989 16 1026 22
<< metal2 >>
rect 109 1254 113 1257
rect 313 1218 407 1221
rect 411 1218 630 1221
rect 313 1217 630 1218
rect 310 1144 622 1146
rect 310 1142 345 1144
rect 350 1142 622 1144
rect 119 1106 130 1110
rect 312 1062 611 1064
rect 312 1060 364 1062
rect 369 1060 611 1062
rect 305 1027 324 1030
rect 321 919 324 1027
rect 607 935 611 1060
rect 618 944 622 1142
rect 626 953 630 1217
rect 626 949 650 953
rect 618 940 652 944
rect 607 931 652 935
rect 350 891 354 894
rect 629 714 633 784
rect 629 711 694 714
rect 629 710 633 711
<< metal3 >>
rect 103 1258 110 1259
rect 103 1253 104 1258
rect 109 1253 110 1258
rect 103 1249 110 1253
rect 104 1112 110 1249
rect 344 1144 351 1145
rect 344 1140 345 1144
rect 350 1140 351 1144
rect 104 1111 120 1112
rect 104 1106 114 1111
rect 119 1106 120 1111
rect 104 1105 120 1106
rect 344 1016 351 1140
rect 295 1010 351 1016
rect 363 1062 370 1063
rect 363 1057 364 1062
rect 369 1057 370 1062
rect 295 900 302 1010
rect 363 1005 370 1057
rect 295 899 355 900
rect 295 894 296 899
rect 301 894 349 899
rect 354 894 355 899
rect 295 893 355 894
<< polycontact >>
rect 406 1008 410 1012
<< m2contact >>
rect 113 1254 117 1258
rect 407 1218 411 1222
rect 130 1106 135 1110
rect 301 1027 305 1031
rect 629 784 633 788
<< m3contact >>
rect 104 1253 109 1258
rect 345 1140 350 1144
rect 114 1106 119 1111
rect 364 1057 369 1062
rect 296 894 301 899
rect 349 894 354 899
use decoder  decoder_0
timestamp 1523195521
transform 1 0 90 0 1 1182
box -58 -160 229 80
use 3seg  3seg_0
timestamp 1523195521
transform 1 0 20 0 1 682
box -20 -682 977 331
use dip2  dip2_1
timestamp 1523195521
transform 1 0 1062 0 1 959
box -35 -277 1713 370
use dip2  dip2_0
timestamp 1523195521
transform 1 0 1052 0 1 285
box -35 -277 1713 370
<< labels >>
rlabel metal1 13 1251 13 1251 1 vdd
rlabel metal1 326 1167 326 1168 1 gnd
rlabel metal1 -17 996 -17 997 3 vdd
rlabel metal1 7 768 7 768 1 gnd
rlabel metal2 684 712 684 713 1 s
<< end >>
