* Spice description of iv1v2x2
* Spice driver version 134999461
* Date 17/05/2007 at  9:11:42
* wsclib 0.13um values
.subckt iv1v2x2 a vdd vss z
M01 vdd   a     z     vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M02 vss   a     z     vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
C3  a     vss   0.353f
C2  z     vss   0.615f
.ends
