* Thu Jan 11 13:03:20 CET 2007
.subckt nr2v0x2 a b vdd vss z
*SPICE circuit <nr2v0x2> from XCircuit v3.20

m1 z a vss vss n w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m2 n1 a vdd vdd p w=56u l=2.3636u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m3 z b vss vss n w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m4 z b n1 vdd p w=56u l=2.3636u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
.ends
