* Tue Feb 20 08:57:11 CET 2007
.subckt iv1v7x4 a vdd vss z
*SPICE circuit <iv1v7x4> from XCircuit v3.20

m1 z a vss vss n w=40u l=2.3636u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m2 z a vdd vdd p w=56u l=2.3636u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
.ends
