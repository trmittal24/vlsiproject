* Spice description of iv1v5x2
* Spice driver version 134999461
* Date 17/05/2007 at  9:13:20
* wsclib 0.13um values
.subckt iv1v5x2 a vdd vss z
M01 vdd   a     z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M02 vss   a     z     vss n  L=0.12U  W=0.605U AS=0.160325P AD=0.160325P PS=1.74U   PD=1.74U
C3  a     vss   0.641f
C2  z     vss   0.840f
.ends
