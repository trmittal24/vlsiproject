* Thu Dec 14 09:40:27 CET 2006
.subckt cgi2bv0x3 a b c vdd vss z
*SPICE circuit <cgi2bv0x3> from XCircuit v3.20

m1 bn b vdd vdd p w=64u l=2.3636u ad='64u*5u+12p' as='64u*5u+12p' pd='64u*2+14u' ps='64u*2+14u'
m2 bn b vss vss n w=32u l=2.3636u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m3 n1 bn vdd vdd p w=84u l=2.3636u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m4 n1 a vdd vdd p w=84u l=2.3636u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m5 z c n1 vdd p w=84u l=2.3636u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m6 n2 a vdd vdd p w=84u l=2.3636u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m7 z bn n2 vdd p w=84u l=2.3636u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m8 n3 bn vss vss n w=42u l=2.3636u ad='42u*5u+12p' as='42u*5u+12p' pd='42u*2+14u' ps='42u*2+14u'
m9 n3 a vss vss n w=42u l=2.3636u ad='42u*5u+12p' as='42u*5u+12p' pd='42u*2+14u' ps='42u*2+14u'
m10 n4 a vss vss n w=42u l=2.3636u ad='42u*5u+12p' as='42u*5u+12p' pd='42u*2+14u' ps='42u*2+14u'
m11 z bn n4 vss n w=42u l=2.3636u ad='42u*5u+12p' as='42u*5u+12p' pd='42u*2+14u' ps='42u*2+14u'
m12 z c n3 vss n w=42u l=2.3636u ad='42u*5u+12p' as='42u*5u+12p' pd='42u*2+14u' ps='42u*2+14u'
.ends
