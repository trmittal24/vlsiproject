* Wed Apr 11 08:44:26 CEST 2007
.subckt xor2v0x05 a b vdd vss z
*SPICE circuit <xor2v0x05> from XCircuit v3.4 rev 26

m1 z bn an vdd p w=13u l=2u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m2 bn b vss vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m3 an a vss vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m4 n1 an vss vss n w=9u l=2u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m5 z bn n1 vss n w=9u l=2u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m6 an a vdd vdd p w=13u l=2u ad='13u*5u+12p' as='13u*5u+12p' pd='13u*2+14u' ps='13u*2+14u'
m7 bn b vdd vdd p w=21u l=2u ad='21u*5u+12p' as='21u*5u+12p' pd='21u*2+14u' ps='21u*2+14u'
m8 z b an vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m9 z an bn vdd p w=21u l=2u ad='21u*5u+12p' as='21u*5u+12p' pd='21u*2+14u' ps='21u*2+14u'
.ends
