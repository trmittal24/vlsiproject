* Wed May  2 18:19:56 CEST 2007
.subckt xnr2v6x1 a b vdd vss z
*SPICE circuit <xnr2v6x1> from XCircuit v3.4 rev 26

m1 an a vdd vdd p w=11u l=2u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m2 an a vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m3 bn b vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m4 bn b vdd vdd p w=11u l=2u ad='11u*5u+12p' as='11u*5u+12p' pd='11u*2+14u' ps='11u*2+14u'
m5 z a n2 vss n w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m6 z an n1 vdd p w=27u l=2u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
m7 n1 a vdd vdd p w=27u l=2u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
m8 n1 bn vdd vdd p w=27u l=2u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
m9 n2 an vss vss n w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m10 n2 bn vss vss n w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m11 z b n2 vss n w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m12 z b n1 vdd p w=27u l=2u ad='27u*5u+12p' as='27u*5u+12p' pd='27u*2+14u' ps='27u*2+14u'
.ends
