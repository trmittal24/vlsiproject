magic
tech scmos
timestamp 1523182099
<< polysilicon >>
rect 152 -101 154 -58
rect 412 -102 414 -59
rect 672 -102 674 -60
<< metal1 >>
rect 60 317 273 320
rect 60 313 130 317
rect 134 313 273 317
rect 60 311 273 313
rect 152 -32 769 -29
rect 152 -54 155 -32
rect 412 -45 753 -42
rect 412 -55 415 -45
rect 676 -60 743 -57
rect -17 -91 16 -88
rect -12 -96 16 -91
rect 217 -156 233 -152
rect 237 -156 240 -152
rect -19 -528 27 -526
rect -19 -533 -8 -528
rect -3 -533 27 -528
rect -19 -534 27 -533
rect 294 -673 334 -670
rect 294 -678 295 -673
rect 300 -678 334 -673
<< metal2 >>
rect 134 313 145 317
rect 733 282 772 286
rect 225 238 233 241
rect 739 199 756 202
rect 733 120 746 123
rect 743 -56 746 120
rect 753 -41 756 199
rect 769 -28 772 282
rect -17 -91 -9 -90
rect -12 -96 -9 -91
rect 233 -152 237 -146
rect 144 -452 150 -449
rect -11 -528 -5 -527
rect -11 -533 -8 -528
rect -16 -534 -5 -533
rect 158 -596 160 -594
rect 164 -596 165 -594
rect 158 -607 165 -596
rect 295 -673 300 -666
<< metal3 >>
rect 144 318 152 319
rect 144 312 145 318
rect 151 312 152 318
rect -18 40 -10 41
rect 144 40 152 312
rect -18 33 152 40
rect -18 -81 -10 33
rect 144 32 152 33
rect 231 242 240 243
rect 231 236 233 242
rect 239 236 240 242
rect 231 235 240 236
rect -18 -82 -8 -81
rect -18 -90 -17 -82
rect -9 -90 -8 -82
rect -18 -91 -8 -90
rect -18 -349 -10 -91
rect -19 -351 -10 -349
rect 231 -140 239 235
rect 231 -146 232 -140
rect 238 -146 239 -140
rect -19 -525 -11 -351
rect 231 -384 239 -146
rect 150 -392 239 -384
rect 150 -438 158 -392
rect 231 -394 239 -392
rect 150 -444 159 -438
rect 149 -446 159 -444
rect 149 -453 150 -446
rect 158 -453 159 -446
rect 149 -454 159 -453
rect -20 -526 -10 -525
rect -20 -533 -19 -526
rect -11 -533 -10 -526
rect -20 -534 -10 -533
rect -19 -606 -11 -534
rect -20 -639 -11 -606
rect 150 -603 159 -454
rect 150 -608 151 -603
rect 158 -608 159 -603
rect 150 -609 159 -608
rect -20 -658 -12 -639
rect -20 -659 22 -658
rect -20 -660 303 -659
rect -20 -666 294 -660
rect 301 -666 303 -660
rect -20 -667 303 -666
<< polycontact >>
rect 152 -58 156 -54
rect 412 -59 416 -55
rect 672 -60 676 -56
<< m2contact >>
rect 130 313 134 317
rect 221 238 225 242
rect 735 198 739 202
rect 769 -32 773 -28
rect 753 -45 757 -41
rect 743 -60 747 -56
rect -17 -96 -12 -91
rect 233 -156 237 -152
rect 140 -452 144 -448
rect -8 -533 -3 -528
rect 160 -596 164 -592
rect 295 -678 300 -673
<< m3contact >>
rect 145 312 151 318
rect 233 236 239 242
rect -17 -90 -9 -82
rect 232 -146 238 -140
rect 150 -453 158 -446
rect -19 -533 -11 -526
rect 151 -608 158 -603
rect 294 -666 301 -660
use firseg  firseg_0
timestamp 1523182099
transform 1 0 0 0 1 80
box 0 -80 739 251
use 2seg  2seg_0
timestamp 1523182099
transform 1 0 2 0 1 -363
box 0 -319 975 298
<< end >>
