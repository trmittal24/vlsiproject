* Spice description of noa3ao322_x4
* Spice driver version 134999461
* Date 21/07/2007 at 19:31:16
* sxlib 0.13um values
.subckt noa3ao322_x4 i0 i1 i2 i3 i4 i5 i6 nq vdd vss
Mtr_00001 vss   sig4  nq    vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00002 nq    sig4  vss   vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00003 sig4  sig8  vss   vss n  L=0.12U  W=0.76U  AS=0.2014P   AD=0.2014P   PS=2.05U   PD=2.05U
Mtr_00004 vss   i5    sig10 vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00005 vss   i3    sig10 vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00006 sig2  i0    vss   vss n  L=0.12U  W=0.87U  AS=0.23055P  AD=0.23055P  PS=2.27U   PD=2.27U
Mtr_00007 sig8  i2    sig9  vss n  L=0.12U  W=0.87U  AS=0.23055P  AD=0.23055P  PS=2.27U   PD=2.27U
Mtr_00008 sig10 i4    vss   vss n  L=0.12U  W=0.43U  AS=0.11395P  AD=0.11395P  PS=1.39U   PD=1.39U
Mtr_00009 sig9  i1    sig2  vss n  L=0.12U  W=0.87U  AS=0.23055P  AD=0.23055P  PS=2.27U   PD=2.27U
Mtr_00010 sig10 i6    sig8  vss n  L=0.12U  W=0.65U  AS=0.17225P  AD=0.17225P  PS=1.83U   PD=1.83U
Mtr_00011 vdd   sig8  sig4  vdd p  L=0.12U  W=1.31U  AS=0.34715P  AD=0.34715P  PS=3.15U   PD=3.15U
Mtr_00012 vdd   i1    sig11 vdd p  L=0.12U  W=1.2U   AS=0.318P    AD=0.318P    PS=2.93U   PD=2.93U
Mtr_00013 sig11 i5    sig13 vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00014 sig13 i4    sig12 vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00015 sig11 i0    vdd   vdd p  L=0.12U  W=1.2U   AS=0.318P    AD=0.318P    PS=2.93U   PD=2.93U
Mtr_00016 nq    sig4  vdd   vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00017 sig11 i2    vdd   vdd p  L=0.12U  W=1.2U   AS=0.318P    AD=0.318P    PS=2.93U   PD=2.93U
Mtr_00018 sig8  i6    sig11 vdd p  L=0.12U  W=1.31U  AS=0.34715P  AD=0.34715P  PS=3.15U   PD=3.15U
Mtr_00019 vdd   sig4  nq    vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00020 sig12 i3    sig8  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
C6  i0    vss   0.676f
C7  i1    vss   0.661f
C18 i2    vss   0.550f
C15 i3    vss   0.676f
C17 i4    vss   0.668f
C16 i5    vss   0.661f
C14 i6    vss   0.592f
C3  nq    vss   0.871f
C10 sig10 vss   0.219f
C11 sig11 vss   0.501f
C4  sig4  vss   0.851f
C8  sig8  vss   1.107f
.ends
