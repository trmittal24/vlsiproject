* Tue Feb 20 08:57:11 CET 2007
.subckt iv1v0x12 a vdd vss z
*SPICE circuit <iv1v0x12> from XCircuit v3.4 rev 26

m1 z a vss vss n w=108u l=2.3636u ad='108u*5u+12p' as='108u*5u+12p' pd='108u*2+14u' ps='108u*2+14u'
m2 z a vdd vdd p w=152u l=2.3636u ad='152u*5u+12p' as='152u*5u+12p' pd='152u*2+14u' ps='152u*2+14u'
.ends
