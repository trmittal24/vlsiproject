* Sat Aug 27 22:10:07 CEST 2005
.subckt iv1v4x6 a vdd vss z 
*SPICE circuit <iv1v4x6> from XCircuit v3.20

m1 z a vss vss n w=24u l=2.3636u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m2 z a vdd vdd p w=96u l=2.3636u ad='96u*5u+12p' as='96u*5u+12p' pd='96u*2+14u' ps='96u*2+14u'
.ends
