* Spice description of or2_x1
* Spice driver version 134999461
* Date 31/05/2007 at 21:35:35
* vxlib 0.13um values
.subckt or2_x1 a b vdd vss z
M1a sig4  a     vdd   vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M1b sig2  b     sig4  vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M1z vdd   sig2  z     vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M2a vss   a     sig2  vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M2b sig2  b     vss   vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M2z z     sig2  vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
C6  a     vss   0.537f
C7  b     vss   0.545f
C2  sig2  vss   0.862f
C3  z     vss   0.872f
.ends
