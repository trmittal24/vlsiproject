* Sat Aug 27 19:28:19 CEST 2005
.subckt nd2v5x1 a b vdd vss z 
*SPICE circuit <nd2v5x1> from XCircuit v3.20

m1 n1 a vss vss n w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m2 z a vdd vdd p w=19u l=2.3636u ad='19u*5u+12p' as='19u*5u+12p' pd='19u*2+14u' ps='19u*2+14u'
m3 z b n1 vss n w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m4 z b vdd vdd p w=19u l=2.3636u ad='19u*5u+12p' as='19u*5u+12p' pd='19u*2+14u' ps='19u*2+14u'
.ends
