* Sat Apr  9 12:32:19 CEST 2005
.subckt or2v0x3 a b vdd vss z 
*SPICE circuit <or2v0x3> from XCircuit v3.20

m1 z zn vdd vdd p w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m2 z zn vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m3 zn a vss vss n w=10u l=2u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m4 n1 a vdd vdd p w=36u l=2u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
m5 zn b vss vss n w=10u l=2u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m6 zn b n1 vdd p w=36u l=2u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
.ends
