* Fri Apr  8 11:37:35 CEST 2005
.subckt aon21bv0x3 a1 a2 b vdd vss z 
*SPICE circuit <aon21bv0x3> from XCircuit v3.20

m1 an a1 vdd vdd p w=25u l=2u ad='25u*5u+12p' as='25u*5u+12p' pd='25u*2+14u' ps='25u*2+14u'
m2 z an vdd vdd p w=34u l=2u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
m3 an a2 vdd vdd p w=25u l=2u ad='25u*5u+12p' as='25u*5u+12p' pd='25u*2+14u' ps='25u*2+14u'
m4 n1 a1 vss vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m5 an a2 n1 vss n w=20u l=2u ad='20u*5u+12p' as='20u*5u+12p' pd='20u*2+14u' ps='20u*2+14u'
m6 z b n2 vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m7 n2 an vss vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m8 z b vdd vdd p w=34u l=2u ad='34u*5u+12p' as='34u*5u+12p' pd='34u*2+14u' ps='34u*2+14u'
.ends
