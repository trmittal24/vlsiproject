* Sat Aug 27 22:10:19 CEST 2005
.subckt iv1v5x6 a vdd vss z 
*SPICE circuit <iv1v5x6> from XCircuit v3.20

m1 z a vss vss n w=32u l=2.3636u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m2 z a vdd vdd p w=84u l=2.3636u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
.ends
