* Spice description of bf1_x4
* Spice driver version 134999461
* Date 31/05/2007 at 21:33:06
* vxlib 0.13um values
.subckt bf1_x4 a vdd vss z
M1a sig3  a     vdd   vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M1b vss   a     sig3  vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
M1z vdd   sig3  z     vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M2z z     sig3  vdd   vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M3z z     sig3  vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
M4z vss   sig3  z     vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
C5  a     vss   0.568f
C3  sig3  vss   0.841f
C2  z     vss   0.923f
.ends
