* Sat Aug 27 22:10:14 CEST 2005
.subckt iv1v5x12 a vdd vss z 
*SPICE circuit <iv1v5x12> from XCircuit v3.20

m1 z a vss vss n w=62u l=2.3636u ad='62u*5u+12p' as='62u*5u+12p' pd='62u*2+14u' ps='62u*2+14u'
m2 z a vdd vdd p w=160u l=2.3636u ad='160u*5u+12p' as='160u*5u+12p' pd='160u*2+14u' ps='160u*2+14u'
.ends
