* Sun Mar 25 12:05:40 CEST 2007
.subckt mxi2v2x05 a0 a1 s vdd vss z
*SPICE circuit <mxi2v2x05> from XCircuit v3.4 rev 26

m1 a0n a0 vdd vdd p w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m2 a1n a1 vdd vdd p w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m3 z sn a1n vdd p w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m4 a0n s z vdd p w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m5 sn s vdd vdd p w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m6 a1n a1 vss vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m7 z sn a0n vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m8 a1n s z vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m9 a0n a0 vss vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m10 sn s vss vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
.ends
