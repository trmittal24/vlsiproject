* Tue Aug 10 11:21:07 CEST 2004
.subckt iv1_x05 a vdd vss z 
*SPICE circuit <iv1_x05> from XCircuit v3.10

m1 z a vss vss n w=6u l=2u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m2 z a vdd vdd p w=12u l=2u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
.ends
