* Tue Aug 10 11:21:07 CEST 2004
.subckt oan22_x2 a1 a2 b1 b2 vdd vss z 
*SPICE circuit <oan22_x2> from XCircuit v3.10

m1 z zn vss vss n w=19u l=2.3636u ad='19u*5u+12p' as='19u*5u+12p' pd='19u*2+14u' ps='19u*2+14u'
m2 z zn vdd vdd p w=39u l=2.3636u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m3 zn b1 n3 vss n w=17u l=2.3636u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m4 n2 b1 vdd vdd p w=39u l=2.3636u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m5 n1 a1 vdd vdd p w=39u l=2.3636u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m6 zn b2 n2 vdd p w=39u l=2.3636u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m7 n3 a2 vss vss n w=17u l=2.3636u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m8 n3 a1 vss vss n w=17u l=2.3636u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m9 zn b2 n3 vss n w=17u l=2.3636u ad='17u*5u+12p' as='17u*5u+12p' pd='17u*2+14u' ps='17u*2+14u'
m10 zn a2 n1 vdd p w=39u l=2.3636u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
.ends
