* Mon Aug 16 14:10:57 CEST 2004
.subckt cgi2v0x05 a b c vdd vss z 
*SPICE circuit <cgi2v0x05> from XCircuit v3.10

m1 n1 b vdd vdd p w=16u l=2u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m2 n2 a vdd vdd p w=16u l=2u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m3 z b n2 vdd p w=16u l=2u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m4 n4 a vss vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m5 z b n4 vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m6 z c n1 vdd p w=16u l=2u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m7 n1 a vdd vdd p w=16u l=2u ad='16u*5u+12p' as='16u*5u+12p' pd='16u*2+14u' ps='16u*2+14u'
m8 n3 b vss vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m9 n3 a vss vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
m10 z c n3 vss n w=7u l=2u ad='7u*5u+12p' as='7u*5u+12p' pd='7u*2+14u' ps='7u*2+14u'
.ends
