* Mon Aug 16 14:10:59 CEST 2004
.subckt nd2v0x1 a b vdd vss z 
*SPICE circuit <nd2v0x1> from XCircuit v3.10

m1 n1 a vss vss n w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m2 z a vdd vdd p w=14u l=2.3636u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m3 z b n1 vss n w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m4 z b vdd vdd p w=14u l=2.3636u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
.ends
