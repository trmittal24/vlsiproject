* Tue Aug 10 11:21:07 CEST 2004
.subckt oai21_x05 a1 a2 b vdd vss z 
*SPICE circuit <oai21_x05> from XCircuit v3.10

m1 n1 a1 vdd vdd p w=23u l=2.3636u ad='23u*5u+12p' as='23u*5u+12p' pd='23u*2+14u' ps='23u*2+14u'
m2 z b vdd vdd p w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m3 n2 a2 vss vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m4 n2 a1 vss vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m5 z b n2 vss n w=10u l=2.3636u ad='10u*5u+12p' as='10u*5u+12p' pd='10u*2+14u' ps='10u*2+14u'
m6 z a2 n1 vdd p w=23u l=2.3636u ad='23u*5u+12p' as='23u*5u+12p' pd='23u*2+14u' ps='23u*2+14u'
.ends
