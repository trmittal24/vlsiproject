* Spice description of oai22_x05
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:10
*
.subckt oai22_x05 a1 a2 b1 b2 vdd vss z 
M1  n1    a1    vdd   vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M2  z     a2    n1    vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M4  n2    b2    z     vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M3  vdd   b1    n2    vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M6  vss   a2    sig1  vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M5  sig1  a1    vss   vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M8  sig1  b2    z     vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
M7  z     b1    sig1  vss n  L=0.13U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U  
C10 a1    vss   1.579f
C9  a2    vss   1.033f
C8  b2    vss   1.343f
C7  b1    vss   1.334f
C4  vdd   vss   1.346f
C2  z     vss   2.763f
C1  sig1  vss   1.266f
.ends
