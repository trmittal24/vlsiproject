magic
tech scmos
timestamp 1520662567
<< pwell >>
rect -66 12 -10 36
rect 0 12 152 36
rect -66 0 152 12
rect -66 -28 14 0
<< nwell >>
rect -66 60 152 80
rect -66 36 -10 60
rect 0 36 152 60
rect -66 -72 14 -28
<< polysilicon >>
rect -52 66 -50 71
rect -42 66 -40 71
rect 13 70 15 74
rect -30 60 -28 65
rect 59 72 115 74
rect 59 64 61 72
rect 69 64 71 68
rect 79 64 81 68
rect 86 64 88 72
rect 96 64 98 68
rect 103 64 105 68
rect 23 56 25 61
rect 42 58 44 63
rect 49 58 51 63
rect -52 38 -50 42
rect -42 38 -40 42
rect -30 39 -28 42
rect -30 38 -23 39
rect -53 32 -47 38
rect -43 37 -37 38
rect -43 33 -42 37
rect -38 33 -37 37
rect -30 34 -28 38
rect -24 34 -23 38
rect -30 33 -23 34
rect 13 38 15 42
rect 23 39 25 42
rect 23 38 38 39
rect 13 37 19 38
rect 23 37 33 38
rect 13 33 14 37
rect 18 33 19 37
rect -43 32 -37 33
rect -50 29 -48 32
rect -43 29 -41 32
rect -29 29 -27 33
rect 13 32 19 33
rect 31 34 33 37
rect 37 34 38 38
rect 31 33 38 34
rect 13 28 15 32
rect 31 30 33 33
rect -29 15 -27 20
rect 42 23 44 52
rect 49 48 51 52
rect 49 47 55 48
rect 49 43 50 47
rect 54 43 55 47
rect 49 42 55 43
rect 59 38 61 52
rect 49 36 61 38
rect 49 23 51 36
rect 69 33 71 52
rect 79 48 81 58
rect 75 47 81 48
rect 75 43 76 47
rect 80 43 81 47
rect 75 42 81 43
rect 69 32 75 33
rect 55 31 61 32
rect 55 27 56 31
rect 60 27 61 31
rect 55 26 61 27
rect 59 23 61 26
rect 69 28 70 32
rect 74 28 75 32
rect 69 27 75 28
rect 69 23 71 27
rect 79 23 81 42
rect 86 38 88 58
rect 113 62 115 72
rect 133 63 135 68
rect 96 48 98 51
rect 92 47 98 48
rect 92 43 93 47
rect 97 43 98 47
rect 92 42 98 43
rect 103 39 105 51
rect 113 48 115 51
rect 133 49 135 53
rect 126 48 135 49
rect 113 46 121 48
rect 119 39 121 46
rect 126 44 127 48
rect 131 44 135 48
rect 126 43 135 44
rect 103 38 109 39
rect 86 36 98 38
rect 86 31 92 32
rect 86 27 87 31
rect 91 27 92 31
rect 86 26 92 27
rect 86 23 88 26
rect 96 23 98 36
rect 103 34 104 38
rect 108 34 109 38
rect 103 33 109 34
rect 119 38 125 39
rect 119 34 120 38
rect 124 34 125 38
rect 119 33 125 34
rect 103 23 105 33
rect 123 30 125 33
rect 133 30 135 43
rect 31 18 33 23
rect 123 19 125 24
rect 133 18 135 23
rect -50 6 -48 10
rect -43 6 -41 10
rect 13 11 15 14
rect 42 11 44 17
rect 49 12 51 17
rect 13 9 44 11
rect 59 8 61 17
rect 69 12 71 17
rect 79 12 81 17
rect 86 8 88 17
rect 96 12 98 17
rect 103 12 105 17
rect 59 6 88 8
rect -51 -2 -49 2
rect -44 -2 -42 2
rect -11 -2 -9 2
rect -4 -2 -2 2
rect -51 -29 -49 -22
rect -44 -25 -42 -22
rect -60 -30 -49 -29
rect -60 -34 -59 -30
rect -55 -34 -49 -30
rect -45 -26 -39 -25
rect -45 -30 -44 -26
rect -40 -30 -39 -26
rect -11 -29 -9 -22
rect -4 -25 -2 -22
rect -45 -31 -39 -30
rect -60 -35 -49 -34
rect -51 -38 -49 -35
rect -41 -38 -39 -31
rect -20 -30 -9 -29
rect -20 -34 -19 -30
rect -15 -34 -9 -30
rect -5 -26 1 -25
rect -5 -30 -4 -26
rect 0 -30 1 -26
rect -5 -31 1 -30
rect -20 -35 -9 -34
rect -11 -38 -9 -35
rect -1 -38 1 -31
rect -51 -66 -49 -62
rect -41 -66 -39 -62
rect -11 -66 -9 -62
rect -1 -66 1 -62
<< ndiffusion >>
rect -55 22 -50 29
rect -57 21 -50 22
rect -57 17 -56 21
rect -52 17 -50 21
rect -57 16 -50 17
rect -55 10 -50 16
rect -48 10 -43 29
rect -41 22 -29 29
rect -41 18 -36 22
rect -32 20 -29 22
rect -27 28 -20 29
rect 24 29 31 30
rect -27 24 -25 28
rect -21 24 -20 28
rect -27 23 -20 24
rect 6 27 13 28
rect 6 23 7 27
rect 11 23 13 27
rect -27 20 -22 23
rect 6 22 13 23
rect -32 18 -31 20
rect -41 15 -31 18
rect -41 11 -36 15
rect -32 11 -31 15
rect 8 14 13 22
rect 15 20 20 28
rect 24 25 25 29
rect 29 25 31 29
rect 24 24 31 25
rect 26 23 31 24
rect 33 23 40 30
rect 116 29 123 30
rect 116 25 117 29
rect 121 25 123 29
rect 116 24 123 25
rect 125 29 133 30
rect 125 25 127 29
rect 131 25 133 29
rect 125 24 133 25
rect 15 19 22 20
rect 15 15 17 19
rect 21 15 22 19
rect 35 22 42 23
rect 35 18 36 22
rect 40 18 42 22
rect 35 17 42 18
rect 44 17 49 23
rect 51 22 59 23
rect 51 18 53 22
rect 57 18 59 22
rect 51 17 59 18
rect 61 22 69 23
rect 61 18 63 22
rect 67 18 69 22
rect 61 17 69 18
rect 71 22 79 23
rect 71 18 73 22
rect 77 18 79 22
rect 71 17 79 18
rect 81 17 86 23
rect 88 22 96 23
rect 88 18 90 22
rect 94 18 96 22
rect 88 17 96 18
rect 98 17 103 23
rect 105 22 112 23
rect 105 18 107 22
rect 111 18 112 22
rect 127 23 133 24
rect 135 29 142 30
rect 135 25 137 29
rect 141 25 142 29
rect 135 23 142 25
rect 105 17 112 18
rect 15 14 22 15
rect -41 10 -31 11
rect -60 -3 -51 -2
rect -60 -7 -59 -3
rect -55 -7 -51 -3
rect -60 -10 -51 -7
rect -60 -14 -59 -10
rect -55 -14 -51 -10
rect -60 -22 -51 -14
rect -49 -22 -44 -2
rect -42 -8 -37 -2
rect -20 -3 -11 -2
rect -20 -7 -19 -3
rect -15 -7 -11 -3
rect -42 -9 -35 -8
rect -42 -13 -40 -9
rect -36 -13 -35 -9
rect -42 -14 -35 -13
rect -20 -10 -11 -7
rect -20 -14 -19 -10
rect -15 -14 -11 -10
rect -42 -22 -37 -14
rect -20 -22 -11 -14
rect -9 -22 -4 -2
rect -2 -8 3 -2
rect -2 -9 5 -8
rect -2 -13 0 -9
rect 4 -13 5 -9
rect -2 -14 5 -13
rect -2 -22 3 -14
<< pdiffusion >>
rect -60 64 -52 66
rect -60 60 -59 64
rect -55 60 -52 64
rect -60 42 -52 60
rect -50 63 -42 66
rect -50 59 -48 63
rect -44 59 -42 63
rect -50 42 -42 59
rect -40 64 -32 66
rect -40 60 -37 64
rect -33 60 -32 64
rect -40 42 -30 60
rect -28 56 -23 60
rect 8 56 13 70
rect -28 55 -21 56
rect -28 51 -26 55
rect -22 51 -21 55
rect -28 50 -21 51
rect 6 54 13 56
rect 6 50 7 54
rect 11 50 13 54
rect -28 42 -23 50
rect 6 47 13 50
rect 6 43 7 47
rect 11 43 13 47
rect 6 42 13 43
rect 15 69 22 70
rect 15 65 17 69
rect 21 65 22 69
rect 15 64 22 65
rect 15 56 21 64
rect 54 58 59 64
rect 34 57 42 58
rect 15 55 23 56
rect 15 51 17 55
rect 21 51 23 55
rect 15 42 23 51
rect 25 48 30 56
rect 34 53 35 57
rect 39 53 42 57
rect 34 52 42 53
rect 44 52 49 58
rect 51 57 59 58
rect 51 53 53 57
rect 57 53 59 57
rect 51 52 59 53
rect 61 57 69 64
rect 61 53 63 57
rect 67 53 69 57
rect 61 52 69 53
rect 71 63 79 64
rect 71 59 73 63
rect 77 59 79 63
rect 71 58 79 59
rect 81 58 86 64
rect 88 63 96 64
rect 88 59 90 63
rect 94 59 96 63
rect 88 58 96 59
rect 71 52 77 58
rect 25 47 32 48
rect 25 43 27 47
rect 31 43 32 47
rect 25 42 32 43
rect 91 51 96 58
rect 98 51 103 64
rect 105 62 110 64
rect 126 62 133 63
rect 105 61 113 62
rect 105 57 107 61
rect 111 57 113 61
rect 105 51 113 57
rect 115 57 120 62
rect 126 58 127 62
rect 131 58 133 62
rect 115 56 122 57
rect 115 52 117 56
rect 121 52 122 56
rect 126 53 133 58
rect 135 59 140 63
rect 135 58 142 59
rect 135 54 137 58
rect 141 54 142 58
rect 135 53 142 54
rect 115 51 122 52
rect -59 -50 -51 -38
rect -59 -54 -57 -50
rect -53 -54 -51 -50
rect -59 -57 -51 -54
rect -59 -61 -57 -57
rect -53 -61 -51 -57
rect -59 -62 -51 -61
rect -49 -43 -41 -38
rect -49 -47 -47 -43
rect -43 -47 -41 -43
rect -49 -50 -41 -47
rect -49 -54 -47 -50
rect -43 -54 -41 -50
rect -49 -62 -41 -54
rect -39 -50 -32 -38
rect -39 -54 -37 -50
rect -33 -54 -32 -50
rect -39 -57 -32 -54
rect -39 -61 -37 -57
rect -33 -61 -32 -57
rect -39 -62 -32 -61
rect -19 -50 -11 -38
rect -19 -54 -17 -50
rect -13 -54 -11 -50
rect -19 -57 -11 -54
rect -19 -61 -17 -57
rect -13 -61 -11 -57
rect -19 -62 -11 -61
rect -9 -43 -1 -38
rect -9 -47 -7 -43
rect -3 -47 -1 -43
rect -9 -50 -1 -47
rect -9 -54 -7 -50
rect -3 -54 -1 -50
rect -9 -62 -1 -54
rect 1 -50 8 -38
rect 1 -54 3 -50
rect 7 -54 8 -50
rect 1 -57 8 -54
rect 1 -61 3 -57
rect 7 -61 8 -57
rect 1 -62 8 -61
<< metal1 >>
rect -64 75 150 76
rect -79 72 150 75
rect -79 68 -27 72
rect -23 69 31 72
rect -23 68 17 69
rect -79 -61 -71 68
rect -59 64 -55 68
rect -37 64 -33 68
rect -59 59 -55 60
rect -52 55 -48 63
rect -44 59 -43 63
rect -37 59 -33 60
rect 21 68 31 69
rect 35 68 41 72
rect 45 68 122 72
rect 126 68 150 72
rect 17 55 21 65
rect -60 49 -48 55
rect -44 51 -26 55
rect -22 51 -21 55
rect 6 54 11 55
rect -60 34 -56 49
rect -60 17 -56 30
rect -52 37 -48 39
rect -44 37 -40 51
rect 6 50 7 54
rect 35 57 39 68
rect 73 63 77 68
rect 73 58 77 59
rect 85 59 90 63
rect 94 59 95 63
rect 106 61 112 68
rect 63 57 67 58
rect 35 52 39 53
rect 42 53 53 57
rect 57 53 58 57
rect 17 50 21 51
rect 6 47 11 50
rect -36 41 -24 47
rect -28 38 -24 41
rect -44 33 -42 37
rect -38 33 -32 37
rect -28 33 -24 34
rect 6 43 7 47
rect 11 43 19 46
rect 6 42 19 43
rect 25 43 27 47
rect 31 43 32 47
rect 6 33 10 42
rect 25 37 29 43
rect 42 38 46 53
rect 63 47 67 53
rect 49 43 50 47
rect 13 33 14 37
rect 18 35 29 37
rect 18 33 25 35
rect -52 29 -48 33
rect -36 29 -32 33
rect -52 25 -40 29
rect -36 28 -20 29
rect -36 25 -25 28
rect -52 17 -51 21
rect -44 17 -40 25
rect -26 24 -25 25
rect -21 24 -20 28
rect 6 28 10 29
rect 32 34 33 38
rect 37 34 48 38
rect 25 29 29 31
rect 6 27 11 28
rect 6 23 7 27
rect 25 24 29 25
rect 6 22 11 23
rect 36 22 40 23
rect -37 18 -36 22
rect -32 18 -31 22
rect -37 15 -31 18
rect -37 12 -36 15
rect -64 11 -36 12
rect -32 12 -31 15
rect 17 19 21 20
rect 17 12 21 15
rect 44 22 48 34
rect 54 32 58 47
rect 63 43 76 47
rect 80 43 81 47
rect 54 31 60 32
rect 54 27 56 31
rect 54 26 60 27
rect 63 22 67 43
rect 85 40 89 59
rect 106 57 107 61
rect 111 57 112 61
rect 126 62 132 68
rect 126 58 127 62
rect 131 58 132 62
rect 137 58 141 59
rect 117 56 121 57
rect 80 36 89 40
rect 93 52 117 54
rect 93 50 121 52
rect 93 47 97 50
rect 125 48 131 54
rect 125 46 127 48
rect 80 33 84 36
rect 70 32 84 33
rect 93 32 97 43
rect 101 38 107 46
rect 117 44 127 46
rect 117 42 131 44
rect 137 38 141 54
rect 101 34 104 38
rect 108 34 112 38
rect 119 34 120 38
rect 124 34 141 38
rect 74 28 84 32
rect 70 27 84 28
rect 44 18 53 22
rect 57 18 58 22
rect 36 12 40 18
rect 63 17 67 18
rect 73 22 77 23
rect 80 22 84 27
rect 87 31 97 32
rect 91 30 97 31
rect 91 29 122 30
rect 91 27 117 29
rect 87 26 117 27
rect 116 25 117 26
rect 121 25 122 29
rect 127 29 131 30
rect 80 18 90 22
rect 94 18 95 22
rect 106 18 107 22
rect 111 18 112 22
rect 73 12 77 18
rect 106 12 112 18
rect 127 12 131 25
rect 137 29 141 34
rect 137 24 141 25
rect -32 11 -26 12
rect -64 8 -26 11
rect -22 8 123 12
rect 127 8 134 12
rect 138 8 150 12
rect -64 4 150 8
rect -64 -3 12 4
rect -64 -4 -59 -3
rect -55 -4 -19 -3
rect -59 -10 -55 -7
rect -15 -4 12 -3
rect -41 -13 -40 -9
rect -59 -15 -55 -14
rect -52 -23 -40 -17
rect -60 -29 -56 -28
rect -44 -26 -40 -23
rect -60 -30 -55 -29
rect -60 -34 -59 -30
rect -44 -31 -40 -30
rect -36 -25 -32 -9
rect -19 -10 -15 -7
rect -1 -13 0 -9
rect -19 -15 -15 -14
rect -12 -18 0 -17
rect -21 -22 0 -18
rect -12 -23 0 -22
rect -36 -28 -16 -25
rect -55 -34 -48 -33
rect -60 -39 -48 -34
rect -36 -41 -32 -28
rect -20 -29 -16 -28
rect -4 -26 0 -23
rect -20 -30 -15 -29
rect -20 -34 -19 -30
rect -4 -31 0 -30
rect 4 -33 8 -9
rect -15 -34 -8 -33
rect -20 -39 -8 -34
rect 4 -36 59 -33
rect 4 -41 8 -36
rect -44 -42 -32 -41
rect -4 -42 8 -41
rect -47 -43 -32 -42
rect -43 -47 -32 -43
rect -7 -43 8 -42
rect -3 -47 8 -43
rect -47 -50 -43 -47
rect -7 -50 -3 -47
rect -58 -54 -57 -50
rect -53 -54 -52 -50
rect -58 -57 -52 -54
rect -47 -55 -43 -54
rect -38 -54 -37 -50
rect -33 -54 -32 -50
rect -58 -60 -57 -57
rect -64 -61 -57 -60
rect -53 -60 -52 -57
rect -38 -57 -32 -54
rect -38 -60 -37 -57
rect -53 -61 -37 -60
rect -33 -60 -32 -57
rect -18 -54 -17 -50
rect -13 -54 -12 -50
rect -18 -57 -12 -54
rect -7 -55 -3 -54
rect 2 -54 3 -50
rect 7 -54 8 -50
rect -18 -60 -17 -57
rect -33 -61 -17 -60
rect -13 -60 -12 -57
rect 2 -57 8 -54
rect 2 -60 3 -57
rect -13 -61 3 -60
rect 7 -60 8 -57
rect 7 -61 12 -60
rect -79 -68 12 -61
<< metal2 >>
rect -59 6 -56 30
rect -52 29 6 33
rect 29 31 30 33
rect -52 28 -48 29
rect -59 1 -22 6
rect -25 -18 -22 1
rect -59 -68 -56 -28
rect 25 -68 30 31
rect 59 -39 63 -37
rect 112 -39 116 34
rect 59 -44 116 -39
rect -59 -71 30 -68
<< ntransistor >>
rect -50 10 -48 29
rect -43 10 -41 29
rect -29 20 -27 29
rect 13 14 15 28
rect 31 23 33 30
rect 123 24 125 30
rect 42 17 44 23
rect 49 17 51 23
rect 59 17 61 23
rect 69 17 71 23
rect 79 17 81 23
rect 86 17 88 23
rect 96 17 98 23
rect 103 17 105 23
rect 133 23 135 30
rect -51 -22 -49 -2
rect -44 -22 -42 -2
rect -11 -22 -9 -2
rect -4 -22 -2 -2
<< ptransistor >>
rect -52 42 -50 66
rect -42 42 -40 66
rect -30 42 -28 60
rect 13 42 15 70
rect 23 42 25 56
rect 42 52 44 58
rect 49 52 51 58
rect 59 52 61 64
rect 69 52 71 64
rect 79 58 81 64
rect 86 58 88 64
rect 96 51 98 64
rect 103 51 105 64
rect 113 51 115 62
rect 133 53 135 63
rect -51 -62 -49 -38
rect -41 -62 -39 -38
rect -11 -62 -9 -38
rect -1 -62 1 -38
<< polycontact >>
rect -42 33 -38 37
rect -28 34 -24 38
rect 14 33 18 37
rect 33 34 37 38
rect 50 43 54 47
rect 76 43 80 47
rect 56 27 60 31
rect 70 28 74 32
rect 93 43 97 47
rect 127 44 131 48
rect 87 27 91 31
rect 104 34 108 38
rect 120 34 124 38
rect -59 -34 -55 -30
rect -44 -30 -40 -26
rect -19 -34 -15 -30
rect -4 -30 0 -26
<< ndcontact >>
rect -56 17 -52 21
rect -36 18 -32 22
rect -25 24 -21 28
rect 7 23 11 27
rect -36 11 -32 15
rect 25 25 29 29
rect 117 25 121 29
rect 127 25 131 29
rect 17 15 21 19
rect 36 18 40 22
rect 53 18 57 22
rect 63 18 67 22
rect 73 18 77 22
rect 90 18 94 22
rect 107 18 111 22
rect 137 25 141 29
rect -59 -7 -55 -3
rect -59 -14 -55 -10
rect -19 -7 -15 -3
rect -40 -13 -36 -9
rect -19 -14 -15 -10
rect 0 -13 4 -9
<< pdcontact >>
rect -59 60 -55 64
rect -48 59 -44 63
rect -37 60 -33 64
rect -26 51 -22 55
rect 7 50 11 54
rect 7 43 11 47
rect 17 65 21 69
rect 17 51 21 55
rect 35 53 39 57
rect 53 53 57 57
rect 63 53 67 57
rect 73 59 77 63
rect 90 59 94 63
rect 27 43 31 47
rect 107 57 111 61
rect 127 58 131 62
rect 117 52 121 56
rect 137 54 141 58
rect -57 -54 -53 -50
rect -57 -61 -53 -57
rect -47 -47 -43 -43
rect -47 -54 -43 -50
rect -37 -54 -33 -50
rect -37 -61 -33 -57
rect -17 -54 -13 -50
rect -17 -61 -13 -57
rect -7 -47 -3 -43
rect -7 -54 -3 -50
rect 3 -54 7 -50
rect 3 -61 7 -57
<< m2contact >>
rect -60 30 -56 34
rect -52 33 -48 37
rect 6 29 10 33
rect 25 31 29 35
rect 112 34 116 38
rect -60 -28 -56 -24
rect -25 -22 -21 -18
rect 59 -37 63 -33
<< psubstratepcontact >>
rect -26 8 -22 12
rect 123 8 127 12
rect 134 8 138 12
<< nsubstratencontact >>
rect -27 68 -23 72
rect 31 68 35 72
rect 41 68 45 72
rect 122 68 126 72
<< psubstratepdiff >>
rect -27 12 -21 13
rect -27 8 -26 12
rect -22 8 -21 12
rect -27 7 -21 8
rect 116 12 145 13
rect 116 8 123 12
rect 127 8 134 12
rect 138 8 145 12
rect 116 7 145 8
<< nsubstratendiff >>
rect -28 72 -22 73
rect -28 68 -27 72
rect -23 68 -22 72
rect 26 72 50 73
rect -28 67 -22 68
rect 26 68 31 72
rect 35 68 41 72
rect 45 68 50 72
rect 26 67 50 68
rect 121 72 127 73
rect 121 68 122 72
rect 126 68 127 72
rect 121 67 127 68
<< labels >>
rlabel polycontact 16 35 16 35 6 zn
rlabel polycontact 34 36 34 36 6 n4
rlabel polycontact 58 29 58 29 6 ci
rlabel polycontact 52 45 52 45 6 ci
rlabel polycontact 72 30 72 30 6 n1
rlabel polycontact 89 29 89 29 6 ci
rlabel polycontact 95 45 95 45 6 ci
rlabel polycontact 78 45 78 45 6 n2
rlabel polycontact 122 36 122 36 6 cn
rlabel metal1 21 35 21 35 6 zn
rlabel metal1 8 40 8 40 6 z
rlabel metal1 16 44 16 44 6 z
rlabel metal1 27 35 27 35 6 zn
rlabel metal1 51 20 51 20 6 n4
rlabel polycontact 57 29 57 29 6 ci
rlabel polycontact 53 45 53 45 6 ci
rlabel metal1 50 55 50 55 6 n4
rlabel metal1 76 8 76 8 6 vss
rlabel metal1 77 30 77 30 6 n1
rlabel metal1 72 45 72 45 6 n2
rlabel metal1 65 37 65 37 6 n2
rlabel metal1 76 72 76 72 6 vdd
rlabel metal1 87 20 87 20 6 n1
rlabel metal1 112 36 112 36 6 d
rlabel metal1 104 40 104 40 6 d
rlabel metal1 95 40 95 40 6 ci
rlabel metal1 90 61 90 61 6 n1
rlabel metal1 104 28 104 28 6 ci
rlabel metal1 130 36 130 36 6 cn
rlabel metal1 120 44 120 44 6 cp
rlabel metal1 128 48 128 48 6 cp
rlabel metal1 139 41 139 41 6 cn
rlabel pdcontact 119 53 119 53 6 ci
rlabel metal1 40 36 40 36 6 n4
rlabel metal1 -38 72 -38 72 6 vdd
rlabel metal1 -33 53 -33 53 6 an
rlabel metal1 -46 -64 -46 -64 2 vdd
rlabel metal1 -46 0 -46 0 2 vss
rlabel metal1 -6 0 -6 0 2 vss
rlabel metal1 -6 -64 -6 -64 2 vdd
rlabel metal1 -50 32 -50 32 6 b
rlabel metal1 -38 8 -38 8 6 vss
rlabel metal1 -10 -36 -10 -36 2 a
rlabel polycontact -18 -32 -18 -32 2 a
rlabel metal1 -42 20 -42 20 6 b
rlabel metal1 -26 40 -26 40 1 k
rlabel metal1 -34 44 -34 44 1 k
rlabel polycontact -40 35 -40 35 1 kn
rlabel polycontact -38 35 -38 35 1 kn
rlabel ntransistor -28 27 -28 27 1 kn
rlabel metal1 -42 -24 -42 -24 1 j
rlabel ntransistor -50 -20 -50 -20 1 j
rlabel metal1 -50 -36 -50 -36 1 q'
rlabel polycontact -58 -32 -58 -32 1 q'
rlabel metal1 -42 -44 -42 -44 1 a
rlabel metal1 -34 -28 -34 -28 1 a
rlabel metal1 6 -28 6 -28 1 c
rlabel metal1 -2 -44 -2 -44 1 c
rlabel ptransistor -50 56 -50 56 1 kq
rlabel metal1 -58 36 -58 36 1 kq
rlabel metal1 -2 -24 -2 -24 1 b4
rlabel ntransistor -10 -20 -10 -20 1 b4
<< end >>
