* SPICE3 file created from totdiff.ext - technology: scmos

.include t14y_tsmc_025_level3.txt

M1000 diff2_0_an2v0x05_0_vdd diff2_2_or2v0x05_0_zn diff2_2_or2v0x05_0_z diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=6096p pd=1908u as=72p ps=38u
M1001 diff2_2_or2v0x05_0_a_24_48# diff2_2_an2v0x05_0_z diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=18u l=2u
+  ad=90p pd=46u as=0p ps=0u
M1002 diff2_2_or2v0x05_0_zn diff2_2_or2v0x05_0_b diff2_2_or2v0x05_0_a_24_48# diff2_0_an2v0x05_0_vdd pfet w=18u l=2u
+  ad=102p pd=50u as=0p ps=0u
M1003 diff2_0_an2v0x05_0_vss diff2_2_or2v0x05_0_zn diff2_2_or2v0x05_0_z diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=3042p pd=1254u as=42p ps=26u
M1004 diff2_2_or2v0x05_0_zn diff2_2_an2v0x05_0_z diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1005 diff2_0_an2v0x05_0_vss diff2_2_or2v0x05_0_b diff2_2_or2v0x05_0_zn diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1006 diff2_0_an2v0x05_0_vdd diff2_2_an2v0x05_0_zn diff2_2_an2v0x05_0_z diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1007 diff2_2_an2v0x05_0_zn diff2_2_an2v0x05_0_a diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1008 diff2_0_an2v0x05_0_vdd diff2_1_or2v0x05_0_z diff2_2_an2v0x05_0_zn diff2_0_an2v0x05_0_vdd pfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1009 diff2_0_an2v0x05_0_vss diff2_2_an2v0x05_0_zn diff2_2_an2v0x05_0_z diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1010 diff2_2_an2v0x05_0_a_23_9# diff2_2_an2v0x05_0_a diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=9u l=2u
+  ad=45p pd=28u as=0p ps=0u
M1011 diff2_2_an2v0x05_0_zn diff2_1_or2v0x05_0_z diff2_2_an2v0x05_0_a_23_9# diff2_0_an2v0x05_0_vss nfet w=9u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1012 diff2_0_an2v0x05_0_vdd diff2_2_xnr2v0x05_0_b diff2_2_xnr2v0x05_0_bn diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1013 diff2_2_xnr2v0x05_0_an diff2_2_an2v0x05_1_b diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1014 diff2_2_an2v0x05_0_a diff2_2_xnr2v0x05_0_b diff2_2_xnr2v0x05_0_an diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=126p pd=52u as=0p ps=0u
M1015 diff2_2_xnr2v0x05_0_a_44_47# diff2_2_xnr2v0x05_0_bn diff2_2_an2v0x05_0_a diff2_0_an2v0x05_0_vdd pfet w=18u l=2u
+  ad=90p pd=46u as=0p ps=0u
M1016 diff2_0_an2v0x05_0_vdd diff2_2_xnr2v0x05_0_an diff2_2_xnr2v0x05_0_a_44_47# diff2_0_an2v0x05_0_vdd pfet w=18u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1017 diff2_0_an2v0x05_0_vss diff2_2_xnr2v0x05_0_b diff2_2_xnr2v0x05_0_bn diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=90p ps=54u
M1018 diff2_2_xnr2v0x05_0_an diff2_2_an2v0x05_1_b diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1019 diff2_2_an2v0x05_0_a diff2_2_xnr2v0x05_0_bn diff2_2_xnr2v0x05_0_an diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1020 diff2_2_xnr2v0x05_0_bn diff2_2_xnr2v0x05_0_an diff2_2_an2v0x05_0_a diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1021 diff2_0_an2v0x05_0_vdd diff2_2_an2v0x05_1_zn diff2_2_or2v0x05_0_b diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1022 diff2_2_an2v0x05_1_zn diff2_2_an2v0x05_1_a diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1023 diff2_0_an2v0x05_0_vdd diff2_2_an2v0x05_1_b diff2_2_an2v0x05_1_zn diff2_0_an2v0x05_0_vdd pfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1024 diff2_0_an2v0x05_0_vss diff2_2_an2v0x05_1_zn diff2_2_or2v0x05_0_b diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1025 diff2_2_an2v0x05_1_a_23_9# diff2_2_an2v0x05_1_a diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=9u l=2u
+  ad=45p pd=28u as=0p ps=0u
M1026 diff2_2_an2v0x05_1_zn diff2_2_an2v0x05_1_b diff2_2_an2v0x05_1_a_23_9# diff2_0_an2v0x05_0_vss nfet w=9u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1027 diff2_2_xor3v0x05_0_a_13_38# diff2_2_an2v0x05_1_a diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=168p pd=68u as=0p ps=0u
M1028 diff2_2_xor3v0x05_0_a_21_38# diff2_2_an2v0x05_1_b diff2_2_xor3v0x05_0_a_13_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=168p pd=68u as=0p ps=0u
M1029 diff2_2_xor3v0x05_0_z diff2_1_or2v0x05_0_z diff2_2_xor3v0x05_0_a_21_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=448p pd=144u as=0p ps=0u
M1030 diff2_2_xor3v0x05_0_a_39_38# diff2_1_or2v0x05_0_z diff2_2_xor3v0x05_0_z diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=140p pd=66u as=0p ps=0u
M1031 diff2_2_an2v0x05_1_a diff2_2_xor3v0x05_0_bn diff2_2_xor3v0x05_0_a_39_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1032 diff2_0_an2v0x05_0_vdd diff2_2_xnr2v0x05_0_b diff2_2_an2v0x05_1_a diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1033 diff2_2_xor3v0x05_0_cn diff2_1_or2v0x05_0_z diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=152p pd=70u as=0p ps=0u
M1034 diff2_2_xor3v0x05_0_bn diff2_2_an2v0x05_1_b diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1035 diff2_2_xor3v0x05_0_a_116_38# diff2_2_xnr2v0x05_0_b diff2_2_xor3v0x05_0_bn diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=140p pd=66u as=0p ps=0u
M1036 diff2_2_xor3v0x05_0_z diff2_2_xor3v0x05_0_cn diff2_2_xor3v0x05_0_a_116_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1037 diff2_2_xor3v0x05_0_a_133_38# diff2_2_xor3v0x05_0_cn diff2_2_xor3v0x05_0_z diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=168p pd=68u as=0p ps=0u
M1038 diff2_2_xor3v0x05_0_a_141_38# diff2_2_xor3v0x05_0_bn diff2_2_xor3v0x05_0_a_133_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=168p pd=68u as=0p ps=0u
M1039 diff2_0_an2v0x05_0_vdd diff2_2_an2v0x05_1_a diff2_2_xor3v0x05_0_a_141_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1040 diff2_2_xor3v0x05_0_a_13_12# diff2_2_an2v0x05_1_a diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=84p pd=40u as=0p ps=0u
M1041 diff2_2_xor3v0x05_0_a_21_12# diff2_2_an2v0x05_1_b diff2_2_xor3v0x05_0_a_13_12# diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=84p pd=40u as=0p ps=0u
M1042 diff2_2_xor3v0x05_0_z diff2_1_or2v0x05_0_z diff2_2_xor3v0x05_0_a_21_12# diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=216p pd=86u as=0p ps=0u
M1043 diff2_2_xor3v0x05_0_a_39_12# diff2_1_or2v0x05_0_z diff2_2_xor3v0x05_0_z diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=109p pd=52u as=0p ps=0u
M1044 diff2_2_an2v0x05_1_a diff2_2_xor3v0x05_0_bn diff2_2_xor3v0x05_0_a_39_12# diff2_0_an2v0x05_0_vss nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1045 diff2_0_an2v0x05_0_vss diff2_2_xnr2v0x05_0_b diff2_2_an2v0x05_1_a diff2_0_an2v0x05_0_vss nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1046 diff2_2_xor3v0x05_0_cn diff2_1_or2v0x05_0_z diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=82p pd=42u as=0p ps=0u
M1047 diff2_2_xor3v0x05_0_bn diff2_2_an2v0x05_1_b diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1048 diff2_2_xor3v0x05_0_a_116_12# diff2_2_xnr2v0x05_0_b diff2_2_xor3v0x05_0_bn diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1049 diff2_2_xor3v0x05_0_z diff2_2_xor3v0x05_0_cn diff2_2_xor3v0x05_0_a_116_12# diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1050 diff2_2_xor3v0x05_0_a_133_12# diff2_2_xor3v0x05_0_cn diff2_2_xor3v0x05_0_z diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=78p pd=38u as=0p ps=0u
M1051 diff2_2_xor3v0x05_0_a_141_12# diff2_2_xor3v0x05_0_bn diff2_2_xor3v0x05_0_a_133_12# diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=78p pd=38u as=0p ps=0u
M1052 diff2_0_an2v0x05_0_vss diff2_2_an2v0x05_1_a diff2_2_xor3v0x05_0_a_141_12# diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1053 diff2_0_an2v0x05_0_vdd diff2_1_or2v0x05_0_zn diff2_1_or2v0x05_0_z diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1054 diff2_1_or2v0x05_0_a_24_48# diff2_1_an2v0x05_0_z diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=18u l=2u
+  ad=90p pd=46u as=0p ps=0u
M1055 diff2_1_or2v0x05_0_zn diff2_1_or2v0x05_0_b diff2_1_or2v0x05_0_a_24_48# diff2_0_an2v0x05_0_vdd pfet w=18u l=2u
+  ad=102p pd=50u as=0p ps=0u
M1056 diff2_0_an2v0x05_0_vss diff2_1_or2v0x05_0_zn diff2_1_or2v0x05_0_z diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1057 diff2_1_or2v0x05_0_zn diff2_1_an2v0x05_0_z diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1058 diff2_0_an2v0x05_0_vss diff2_1_or2v0x05_0_b diff2_1_or2v0x05_0_zn diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1059 diff2_0_an2v0x05_0_vdd diff2_1_an2v0x05_0_zn diff2_1_an2v0x05_0_z diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1060 diff2_1_an2v0x05_0_zn diff2_1_an2v0x05_0_a diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1061 diff2_0_an2v0x05_0_vdd diff2_0_or2v0x05_0_z diff2_1_an2v0x05_0_zn diff2_0_an2v0x05_0_vdd pfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1062 diff2_0_an2v0x05_0_vss diff2_1_an2v0x05_0_zn diff2_1_an2v0x05_0_z diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1063 diff2_1_an2v0x05_0_a_23_9# diff2_1_an2v0x05_0_a diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=9u l=2u
+  ad=45p pd=28u as=0p ps=0u
M1064 diff2_1_an2v0x05_0_zn diff2_0_or2v0x05_0_z diff2_1_an2v0x05_0_a_23_9# diff2_0_an2v0x05_0_vss nfet w=9u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1065 diff2_0_an2v0x05_0_vdd diff2_1_xnr2v0x05_0_b diff2_1_xnr2v0x05_0_bn diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1066 diff2_1_xnr2v0x05_0_an diff2_1_an2v0x05_1_b diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1067 diff2_1_an2v0x05_0_a diff2_1_xnr2v0x05_0_b diff2_1_xnr2v0x05_0_an diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=126p pd=52u as=0p ps=0u
M1068 diff2_1_xnr2v0x05_0_a_44_47# diff2_1_xnr2v0x05_0_bn diff2_1_an2v0x05_0_a diff2_0_an2v0x05_0_vdd pfet w=18u l=2u
+  ad=90p pd=46u as=0p ps=0u
M1069 diff2_0_an2v0x05_0_vdd diff2_1_xnr2v0x05_0_an diff2_1_xnr2v0x05_0_a_44_47# diff2_0_an2v0x05_0_vdd pfet w=18u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1070 diff2_0_an2v0x05_0_vss diff2_1_xnr2v0x05_0_b diff2_1_xnr2v0x05_0_bn diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=90p ps=54u
M1071 diff2_1_xnr2v0x05_0_an diff2_1_an2v0x05_1_b diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1072 diff2_1_an2v0x05_0_a diff2_1_xnr2v0x05_0_bn diff2_1_xnr2v0x05_0_an diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1073 diff2_1_xnr2v0x05_0_bn diff2_1_xnr2v0x05_0_an diff2_1_an2v0x05_0_a diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1074 diff2_0_an2v0x05_0_vdd diff2_1_an2v0x05_1_zn diff2_1_or2v0x05_0_b diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1075 diff2_1_an2v0x05_1_zn diff2_1_an2v0x05_1_a diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1076 diff2_0_an2v0x05_0_vdd diff2_1_an2v0x05_1_b diff2_1_an2v0x05_1_zn diff2_0_an2v0x05_0_vdd pfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1077 diff2_0_an2v0x05_0_vss diff2_1_an2v0x05_1_zn diff2_1_or2v0x05_0_b diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1078 diff2_1_an2v0x05_1_a_23_9# diff2_1_an2v0x05_1_a diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=9u l=2u
+  ad=45p pd=28u as=0p ps=0u
M1079 diff2_1_an2v0x05_1_zn diff2_1_an2v0x05_1_b diff2_1_an2v0x05_1_a_23_9# diff2_0_an2v0x05_0_vss nfet w=9u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1080 diff2_1_xor3v0x05_0_a_13_38# diff2_1_an2v0x05_1_a diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=168p pd=68u as=0p ps=0u
M1081 diff2_1_xor3v0x05_0_a_21_38# diff2_1_an2v0x05_1_b diff2_1_xor3v0x05_0_a_13_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=168p pd=68u as=0p ps=0u
M1082 diff2_1_xor3v0x05_0_z diff2_0_or2v0x05_0_z diff2_1_xor3v0x05_0_a_21_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=448p pd=144u as=0p ps=0u
M1083 diff2_1_xor3v0x05_0_a_39_38# diff2_0_or2v0x05_0_z diff2_1_xor3v0x05_0_z diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=140p pd=66u as=0p ps=0u
M1084 diff2_1_an2v0x05_1_a diff2_1_xor3v0x05_0_bn diff2_1_xor3v0x05_0_a_39_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1085 diff2_0_an2v0x05_0_vdd diff2_1_xnr2v0x05_0_b diff2_1_an2v0x05_1_a diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1086 diff2_1_xor3v0x05_0_cn diff2_0_or2v0x05_0_z diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=152p pd=70u as=0p ps=0u
M1087 diff2_1_xor3v0x05_0_bn diff2_1_an2v0x05_1_b diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1088 diff2_1_xor3v0x05_0_a_116_38# diff2_1_xnr2v0x05_0_b diff2_1_xor3v0x05_0_bn diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=140p pd=66u as=0p ps=0u
M1089 diff2_1_xor3v0x05_0_z diff2_1_xor3v0x05_0_cn diff2_1_xor3v0x05_0_a_116_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1090 diff2_1_xor3v0x05_0_a_133_38# diff2_1_xor3v0x05_0_cn diff2_1_xor3v0x05_0_z diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=168p pd=68u as=0p ps=0u
M1091 diff2_1_xor3v0x05_0_a_141_38# diff2_1_xor3v0x05_0_bn diff2_1_xor3v0x05_0_a_133_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=168p pd=68u as=0p ps=0u
M1092 diff2_0_an2v0x05_0_vdd diff2_1_an2v0x05_1_a diff2_1_xor3v0x05_0_a_141_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1093 diff2_1_xor3v0x05_0_a_13_12# diff2_1_an2v0x05_1_a diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=84p pd=40u as=0p ps=0u
M1094 diff2_1_xor3v0x05_0_a_21_12# diff2_1_an2v0x05_1_b diff2_1_xor3v0x05_0_a_13_12# diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=84p pd=40u as=0p ps=0u
M1095 diff2_1_xor3v0x05_0_z diff2_0_or2v0x05_0_z diff2_1_xor3v0x05_0_a_21_12# diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=216p pd=86u as=0p ps=0u
M1096 diff2_1_xor3v0x05_0_a_39_12# diff2_0_or2v0x05_0_z diff2_1_xor3v0x05_0_z diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=109p pd=52u as=0p ps=0u
M1097 diff2_1_an2v0x05_1_a diff2_1_xor3v0x05_0_bn diff2_1_xor3v0x05_0_a_39_12# diff2_0_an2v0x05_0_vss nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1098 diff2_0_an2v0x05_0_vss diff2_1_xnr2v0x05_0_b diff2_1_an2v0x05_1_a diff2_0_an2v0x05_0_vss nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1099 diff2_1_xor3v0x05_0_cn diff2_0_or2v0x05_0_z diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=82p pd=42u as=0p ps=0u
M1100 diff2_1_xor3v0x05_0_bn diff2_1_an2v0x05_1_b diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1101 diff2_1_xor3v0x05_0_a_116_12# diff2_1_xnr2v0x05_0_b diff2_1_xor3v0x05_0_bn diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1102 diff2_1_xor3v0x05_0_z diff2_1_xor3v0x05_0_cn diff2_1_xor3v0x05_0_a_116_12# diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1103 diff2_1_xor3v0x05_0_a_133_12# diff2_1_xor3v0x05_0_cn diff2_1_xor3v0x05_0_z diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=78p pd=38u as=0p ps=0u
M1104 diff2_1_xor3v0x05_0_a_141_12# diff2_1_xor3v0x05_0_bn diff2_1_xor3v0x05_0_a_133_12# diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=78p pd=38u as=0p ps=0u
M1105 diff2_0_an2v0x05_0_vss diff2_1_an2v0x05_1_a diff2_1_xor3v0x05_0_a_141_12# diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1106 diff2_0_an2v0x05_0_vdd diff2_0_or2v0x05_0_zn diff2_0_or2v0x05_0_z diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1107 diff2_0_or2v0x05_0_a_24_48# diff2_0_an2v0x05_0_z diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=18u l=2u
+  ad=90p pd=46u as=0p ps=0u
M1108 diff2_0_or2v0x05_0_zn diff2_0_or2v0x05_0_b diff2_0_or2v0x05_0_a_24_48# diff2_0_an2v0x05_0_vdd pfet w=18u l=2u
+  ad=102p pd=50u as=0p ps=0u
M1109 diff2_0_an2v0x05_0_vss diff2_0_or2v0x05_0_zn diff2_0_or2v0x05_0_z diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1110 diff2_0_or2v0x05_0_zn diff2_0_an2v0x05_0_z diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1111 diff2_0_an2v0x05_0_vss diff2_0_or2v0x05_0_b diff2_0_or2v0x05_0_zn diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1112 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_zn diff2_0_an2v0x05_0_z diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1113 diff2_0_an2v0x05_0_zn diff2_0_an2v0x05_0_a diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1114 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_b diff2_0_an2v0x05_0_zn diff2_0_an2v0x05_0_vdd pfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1115 diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_zn diff2_0_an2v0x05_0_z diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1116 diff2_0_an2v0x05_0_a_23_9# diff2_0_an2v0x05_0_a diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=9u l=2u
+  ad=45p pd=28u as=0p ps=0u
M1117 diff2_0_an2v0x05_0_zn diff2_0_an2v0x05_0_b diff2_0_an2v0x05_0_a_23_9# diff2_0_an2v0x05_0_vss nfet w=9u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1118 diff2_0_an2v0x05_0_vdd diff2_0_xnr2v0x05_0_b diff2_0_xnr2v0x05_0_bn diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1119 diff2_0_xnr2v0x05_0_an diff2_0_an2v0x05_1_b diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1120 diff2_0_an2v0x05_0_a diff2_0_xnr2v0x05_0_b diff2_0_xnr2v0x05_0_an diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=126p pd=52u as=0p ps=0u
M1121 diff2_0_xnr2v0x05_0_a_44_47# diff2_0_xnr2v0x05_0_bn diff2_0_an2v0x05_0_a diff2_0_an2v0x05_0_vdd pfet w=18u l=2u
+  ad=90p pd=46u as=0p ps=0u
M1122 diff2_0_an2v0x05_0_vdd diff2_0_xnr2v0x05_0_an diff2_0_xnr2v0x05_0_a_44_47# diff2_0_an2v0x05_0_vdd pfet w=18u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1123 diff2_0_an2v0x05_0_vss diff2_0_xnr2v0x05_0_b diff2_0_xnr2v0x05_0_bn diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=90p ps=54u
M1124 diff2_0_xnr2v0x05_0_an diff2_0_an2v0x05_1_b diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1125 diff2_0_an2v0x05_0_a diff2_0_xnr2v0x05_0_bn diff2_0_xnr2v0x05_0_an diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1126 diff2_0_xnr2v0x05_0_bn diff2_0_xnr2v0x05_0_an diff2_0_an2v0x05_0_a diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1127 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_1_zn diff2_0_or2v0x05_0_b diff2_0_an2v0x05_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1128 diff2_0_an2v0x05_1_zn diff2_0_an2v0x05_1_a diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1129 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_1_b diff2_0_an2v0x05_1_zn diff2_0_an2v0x05_0_vdd pfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1130 diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_1_zn diff2_0_or2v0x05_0_b diff2_0_an2v0x05_0_vss nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1131 diff2_0_an2v0x05_1_a_23_9# diff2_0_an2v0x05_1_a diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=9u l=2u
+  ad=45p pd=28u as=0p ps=0u
M1132 diff2_0_an2v0x05_1_zn diff2_0_an2v0x05_1_b diff2_0_an2v0x05_1_a_23_9# diff2_0_an2v0x05_0_vss nfet w=9u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1133 diff2_0_xor3v0x05_0_a_13_38# diff2_0_an2v0x05_1_a diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=168p pd=68u as=0p ps=0u
M1134 diff2_0_xor3v0x05_0_a_21_38# diff2_0_an2v0x05_1_b diff2_0_xor3v0x05_0_a_13_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=168p pd=68u as=0p ps=0u
M1135 diff2_0_xor3v0x05_0_z diff2_0_an2v0x05_0_b diff2_0_xor3v0x05_0_a_21_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=448p pd=144u as=0p ps=0u
M1136 diff2_0_xor3v0x05_0_a_39_38# diff2_0_an2v0x05_0_b diff2_0_xor3v0x05_0_z diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=140p pd=66u as=0p ps=0u
M1137 diff2_0_an2v0x05_1_a diff2_0_xor3v0x05_0_bn diff2_0_xor3v0x05_0_a_39_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1138 diff2_0_an2v0x05_0_vdd diff2_0_xnr2v0x05_0_b diff2_0_an2v0x05_1_a diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1139 diff2_0_xor3v0x05_0_cn diff2_0_an2v0x05_0_b diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=152p pd=70u as=0p ps=0u
M1140 diff2_0_xor3v0x05_0_bn diff2_0_an2v0x05_1_b diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1141 diff2_0_xor3v0x05_0_a_116_38# diff2_0_xnr2v0x05_0_b diff2_0_xor3v0x05_0_bn diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=140p pd=66u as=0p ps=0u
M1142 diff2_0_xor3v0x05_0_z diff2_0_xor3v0x05_0_cn diff2_0_xor3v0x05_0_a_116_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1143 diff2_0_xor3v0x05_0_a_133_38# diff2_0_xor3v0x05_0_cn diff2_0_xor3v0x05_0_z diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=168p pd=68u as=0p ps=0u
M1144 diff2_0_xor3v0x05_0_a_141_38# diff2_0_xor3v0x05_0_bn diff2_0_xor3v0x05_0_a_133_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=168p pd=68u as=0p ps=0u
M1145 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_1_a diff2_0_xor3v0x05_0_a_141_38# diff2_0_an2v0x05_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1146 diff2_0_xor3v0x05_0_a_13_12# diff2_0_an2v0x05_1_a diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=84p pd=40u as=0p ps=0u
M1147 diff2_0_xor3v0x05_0_a_21_12# diff2_0_an2v0x05_1_b diff2_0_xor3v0x05_0_a_13_12# diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=84p pd=40u as=0p ps=0u
M1148 diff2_0_xor3v0x05_0_z diff2_0_an2v0x05_0_b diff2_0_xor3v0x05_0_a_21_12# diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=216p pd=86u as=0p ps=0u
M1149 diff2_0_xor3v0x05_0_a_39_12# diff2_0_an2v0x05_0_b diff2_0_xor3v0x05_0_z diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=109p pd=52u as=0p ps=0u
M1150 diff2_0_an2v0x05_1_a diff2_0_xor3v0x05_0_bn diff2_0_xor3v0x05_0_a_39_12# diff2_0_an2v0x05_0_vss nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1151 diff2_0_an2v0x05_0_vss diff2_0_xnr2v0x05_0_b diff2_0_an2v0x05_1_a diff2_0_an2v0x05_0_vss nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1152 diff2_0_xor3v0x05_0_cn diff2_0_an2v0x05_0_b diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=14u l=2u
+  ad=82p pd=42u as=0p ps=0u
M1153 diff2_0_xor3v0x05_0_bn diff2_0_an2v0x05_1_b diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1154 diff2_0_xor3v0x05_0_a_116_12# diff2_0_xnr2v0x05_0_b diff2_0_xor3v0x05_0_bn diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1155 diff2_0_xor3v0x05_0_z diff2_0_xor3v0x05_0_cn diff2_0_xor3v0x05_0_a_116_12# diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1156 diff2_0_xor3v0x05_0_a_133_12# diff2_0_xor3v0x05_0_cn diff2_0_xor3v0x05_0_z diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=78p pd=38u as=0p ps=0u
M1157 diff2_0_xor3v0x05_0_a_141_12# diff2_0_xor3v0x05_0_bn diff2_0_xor3v0x05_0_a_133_12# diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=78p pd=38u as=0p ps=0u
M1158 diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_1_a diff2_0_xor3v0x05_0_a_141_12# diff2_0_an2v0x05_0_vss nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 diff2_2_xor3v0x05_0_a_141_38# diff2_2_an2v0x05_1_a 2.3fF
C1 diff2_0_an2v0x05_0_vss diff2_1_an2v0x05_1_b 30.5fF
C2 diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_z 8.0fF
C3 diff2_0_an2v0x05_0_vdd diff2_2_an2v0x05_1_zn 6.0fF
C4 diff2_0_or2v0x05_0_z diff2_1_xnr2v0x05_0_b 2.5fF
C5 diff2_0_an2v0x05_0_vss diff2_0_xor3v0x05_0_bn 21.9fF
C6 diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_1_a 19.4fF
C7 diff2_0_xnr2v0x05_0_b diff2_0_an2v0x05_0_b 2.5fF
C8 diff2_0_an2v0x05_0_vss diff2_0_xnr2v0x05_0_an 4.2fF
C9 diff2_0_an2v0x05_0_vdd diff2_0_xnr2v0x05_0_b 31.8fF
C10 diff2_0_an2v0x05_0_vss diff2_2_xnr2v0x05_0_an 4.2fF
C11 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_b 18.6fF
C12 diff2_1_an2v0x05_0_z diff2_0_an2v0x05_0_vss 8.0fF
C13 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_a 22.2fF
C14 diff2_0_an2v0x05_0_vss diff2_0_or2v0x05_0_z 40.7fF
C15 diff2_0_an2v0x05_0_vdd diff2_1_an2v0x05_1_a 48.6fF
C16 diff2_0_an2v0x05_0_vdd diff2_1_an2v0x05_0_zn 6.0fF
C17 diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_zn 9.1fF
C18 diff2_1_xor3v0x05_0_cn diff2_1_an2v0x05_1_b 5.8fF
C19 diff2_0_an2v0x05_1_b diff2_0_xor3v0x05_0_bn 4.0fF
C20 diff2_0_an2v0x05_0_vss diff2_1_xor3v0x05_0_bn 21.9fF
C21 diff2_0_an2v0x05_0_vss diff2_2_or2v0x05_0_z 2.5fF
C22 diff2_1_xor3v0x05_0_z diff2_1_an2v0x05_1_b 4.6fF
C23 diff2_0_an2v0x05_0_vdd diff2_2_or2v0x05_0_zn 11.9fF
C24 diff2_0_an2v0x05_1_a diff2_0_an2v0x05_1_b 5.4fF
C25 diff2_0_an2v0x05_0_vdd diff2_2_or2v0x05_0_b 16.5fF
C26 diff2_0_an2v0x05_0_vdd diff2_2_xor3v0x05_0_bn 10.0fF
C27 diff2_0_an2v0x05_0_vdd diff2_2_xnr2v0x05_0_bn 8.3fF
C28 diff2_0_an2v0x05_0_vdd diff2_0_or2v0x05_0_b 16.5fF
C29 diff2_0_an2v0x05_0_vdd diff2_1_or2v0x05_0_zn 11.9fF
C30 diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_1_zn 9.1fF
C31 diff2_2_an2v0x05_0_a diff2_0_an2v0x05_0_vss 8.0fF
C32 diff2_0_an2v0x05_0_vdd diff2_1_xnr2v0x05_0_b 31.8fF
C33 diff2_2_an2v0x05_1_zn diff2_0_an2v0x05_0_vss 9.1fF
C34 diff2_0_an2v0x05_0_vdd diff2_1_an2v0x05_0_a 22.2fF
C35 diff2_0_an2v0x05_0_vdd diff2_0_xor3v0x05_0_z 17.2fF
C36 diff2_0_an2v0x05_0_vdd diff2_2_xnr2v0x05_0_b 31.8fF
C37 diff2_0_an2v0x05_0_b diff2_0_xor3v0x05_0_cn 5.1fF
C38 diff2_0_an2v0x05_0_vdd diff2_2_an2v0x05_1_b 31.9fF
C39 diff2_0_xor3v0x05_0_a_141_38# diff2_0_an2v0x05_1_a 2.3fF
C40 diff2_0_an2v0x05_0_vdd diff2_0_xor3v0x05_0_cn 17.9fF
C41 diff2_0_an2v0x05_0_vss diff2_0_xnr2v0x05_0_b 70.8fF
C42 diff2_0_or2v0x05_0_z diff2_1_xor3v0x05_0_cn 5.1fF
C43 diff2_0_an2v0x05_0_vdd diff2_2_an2v0x05_0_zn 6.0fF
C44 diff2_0_an2v0x05_0_vdd diff2_1_xnr2v0x05_0_an 11.7fF
C45 diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_b 37.2fF
C46 diff2_1_xor3v0x05_0_cn diff2_1_xor3v0x05_0_bn 2.2fF
C47 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_vss 7.4fF
C48 diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_0_a 8.0fF
C49 diff2_2_xnr2v0x05_0_bn diff2_2_xnr2v0x05_0_b 2.1fF
C50 diff2_1_xor3v0x05_0_z diff2_1_xor3v0x05_0_bn 4.1fF
C51 diff2_2_an2v0x05_1_b diff2_2_xor3v0x05_0_bn 4.0fF
C52 diff2_0_an2v0x05_0_vss diff2_1_an2v0x05_1_a 19.4fF
C53 diff2_0_an2v0x05_0_vss diff2_1_an2v0x05_0_zn 9.1fF
C54 diff2_2_an2v0x05_0_z diff2_0_an2v0x05_0_vdd 12.4fF
C55 diff2_0_an2v0x05_0_vdd diff2_2_an2v0x05_1_a 48.6fF
C56 diff2_0_an2v0x05_0_vdd diff2_1_or2v0x05_0_z 48.5fF
C57 diff2_2_or2v0x05_0_zn diff2_0_an2v0x05_0_vss 8.1fF
C58 diff2_0_an2v0x05_0_vdd diff2_2_xor3v0x05_0_cn 17.9fF
C59 diff2_0_an2v0x05_0_vdd diff2_0_or2v0x05_0_zn 11.9fF
C60 diff2_2_or2v0x05_0_b diff2_0_an2v0x05_0_vss 17.6fF
C61 diff2_1_xor3v0x05_0_a_141_38# diff2_1_an2v0x05_1_a 2.3fF
C62 diff2_0_an2v0x05_0_vss diff2_2_xor3v0x05_0_bn 21.9fF
C63 diff2_2_xnr2v0x05_0_bn diff2_0_an2v0x05_0_vss 26.6fF
C64 diff2_0_an2v0x05_0_vss diff2_0_or2v0x05_0_b 16.3fF
C65 diff2_0_or2v0x05_0_z diff2_1_an2v0x05_1_b 6.8fF
C66 diff2_0_an2v0x05_0_vss diff2_1_or2v0x05_0_zn 8.1fF
C67 diff2_0_an2v0x05_0_vss diff2_1_xnr2v0x05_0_b 70.8fF
C68 diff2_0_an2v0x05_1_b diff2_0_an2v0x05_0_b 6.8fF
C69 diff2_0_an2v0x05_0_vdd diff2_1_an2v0x05_1_zn 6.0fF
C70 diff2_0_an2v0x05_0_vss diff2_1_an2v0x05_0_a 8.0fF
C71 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_1_b 31.9fF
C72 diff2_0_an2v0x05_0_vss diff2_0_xor3v0x05_0_z 4.8fF
C73 diff2_1_an2v0x05_1_b diff2_1_xor3v0x05_0_bn 4.0fF
C74 diff2_2_xnr2v0x05_0_b diff2_0_an2v0x05_0_vss 70.8fF
C75 diff2_0_an2v0x05_0_vdd diff2_1_xnr2v0x05_0_bn 8.3fF
C76 diff2_1_or2v0x05_0_z diff2_2_xor3v0x05_0_bn 2.7fF
C77 diff2_0_an2v0x05_0_vdd diff2_2_xor3v0x05_0_z 17.2fF
C78 diff2_2_xor3v0x05_0_cn diff2_2_xor3v0x05_0_bn 2.2fF
C79 diff2_0_an2v0x05_0_vdd diff2_1_xor3v0x05_0_cn 17.9fF
C80 diff2_0_an2v0x05_0_vss diff2_2_an2v0x05_1_b 30.5fF
C81 diff2_0_an2v0x05_0_vss diff2_0_xor3v0x05_0_cn 15.4fF
C82 diff2_0_an2v0x05_0_vdd diff2_1_xor3v0x05_0_z 17.2fF
C83 diff2_2_an2v0x05_0_zn diff2_0_an2v0x05_0_vss 9.1fF
C84 diff2_0_an2v0x05_0_vss diff2_1_xnr2v0x05_0_an 4.2fF
C85 diff2_0_xnr2v0x05_0_bn diff2_0_xnr2v0x05_0_b 2.1fF
C86 diff2_1_an2v0x05_0_z diff2_0_or2v0x05_0_z 2.0fF
C87 diff2_1_xor3v0x05_0_z diff2_1_an2v0x05_1_a 7.8fF
C88 diff2_1_or2v0x05_0_z diff2_2_xnr2v0x05_0_b 2.5fF
C89 diff2_2_an2v0x05_1_a diff2_2_an2v0x05_1_b 5.4fF
C90 diff2_1_or2v0x05_0_z diff2_2_an2v0x05_1_b 6.8fF
C91 diff2_0_an2v0x05_0_vdd diff2_1_or2v0x05_0_b 16.5fF
C92 diff2_2_xor3v0x05_0_cn diff2_2_an2v0x05_1_b 5.8fF
C93 diff2_2_xor3v0x05_0_z diff2_2_xor3v0x05_0_bn 4.1fF
C94 diff2_0_an2v0x05_0_vdd diff2_0_xnr2v0x05_0_bn 8.3fF
C95 diff2_1_or2v0x05_0_z diff2_2_an2v0x05_0_zn 2.7fF
C96 diff2_1_xnr2v0x05_0_bn diff2_1_xnr2v0x05_0_b 2.1fF
C97 diff2_0_or2v0x05_0_z diff2_1_xor3v0x05_0_bn 2.7fF
C98 diff2_2_an2v0x05_0_z diff2_0_an2v0x05_0_vss 8.0fF
C99 diff2_0_an2v0x05_1_b diff2_0_xor3v0x05_0_z 4.6fF
C100 diff2_0_an2v0x05_0_vss diff2_2_an2v0x05_1_a 19.4fF
C101 diff2_1_or2v0x05_0_z diff2_0_an2v0x05_0_vss 42.2fF
C102 diff2_2_xor3v0x05_0_cn diff2_0_an2v0x05_0_vss 15.4fF
C103 diff2_0_an2v0x05_0_vss diff2_0_or2v0x05_0_zn 8.1fF
C104 diff2_0_an2v0x05_0_vdd diff2_1_an2v0x05_1_b 31.9fF
C105 diff2_2_xor3v0x05_0_z diff2_2_an2v0x05_1_b 4.6fF
C106 diff2_0_an2v0x05_1_b diff2_0_xor3v0x05_0_cn 5.8fF
C107 diff2_0_xor3v0x05_0_bn diff2_0_an2v0x05_0_b 2.7fF
C108 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_z 12.4fF
C109 diff2_1_an2v0x05_1_a diff2_1_an2v0x05_1_b 5.4fF
C110 diff2_0_an2v0x05_0_vdd diff2_0_xor3v0x05_0_bn 10.0fF
C111 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_1_a 48.6fF
C112 diff2_0_an2v0x05_0_vdd diff2_0_xnr2v0x05_0_an 11.7fF
C113 diff2_2_xor3v0x05_0_cn diff2_1_or2v0x05_0_z 5.1fF
C114 diff2_0_an2v0x05_0_vss diff2_1_an2v0x05_1_zn 9.1fF
C115 diff2_0_an2v0x05_0_vss diff2_0_an2v0x05_1_b 30.5fF
C116 diff2_1_xnr2v0x05_0_bn diff2_0_an2v0x05_0_vss 26.6fF
C117 diff2_0_an2v0x05_0_vss diff2_2_xor3v0x05_0_z 4.8fF
C118 diff2_0_an2v0x05_0_vss diff2_1_xor3v0x05_0_cn 15.4fF
C119 diff2_0_an2v0x05_0_vdd diff2_2_xnr2v0x05_0_an 11.7fF
C120 diff2_0_an2v0x05_0_vdd diff2_1_an2v0x05_0_z 12.4fF
C121 diff2_0_an2v0x05_0_vss diff2_1_xor3v0x05_0_z 4.8fF
C122 diff2_2_xor3v0x05_0_z diff2_2_an2v0x05_1_a 7.8fF
C123 diff2_0_an2v0x05_0_vdd diff2_0_or2v0x05_0_z 47.7fF
C124 diff2_0_an2v0x05_0_zn diff2_0_an2v0x05_0_b 2.2fF
C125 diff2_0_an2v0x05_0_vss diff2_1_or2v0x05_0_b 17.0fF
C126 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_0_zn 6.0fF
C127 diff2_0_or2v0x05_0_z diff2_1_an2v0x05_0_zn 3.0fF
C128 diff2_0_xnr2v0x05_0_bn diff2_0_an2v0x05_0_vss 26.6fF
C129 diff2_0_xor3v0x05_0_bn diff2_0_xor3v0x05_0_z 4.1fF
C130 diff2_0_an2v0x05_0_vdd diff2_1_xor3v0x05_0_bn 10.0fF
C131 diff2_0_an2v0x05_0_vdd diff2_2_or2v0x05_0_z 4.4fF
C132 diff2_0_an2v0x05_1_a diff2_0_xor3v0x05_0_z 7.8fF
C133 diff2_0_xor3v0x05_0_bn diff2_0_xor3v0x05_0_cn 2.2fF
C134 diff2_0_an2v0x05_0_vdd diff2_0_an2v0x05_1_zn 6.0fF
C135 diff2_0_an2v0x05_0_vdd diff2_2_an2v0x05_0_a 22.2fF
C136 diff2_0_or2v0x05_0_b 0 2.9fF
C137 diff2_1_or2v0x05_0_b 0 2.9fF
C138 diff2_1_or2v0x05_0_z 0 7.7fF
C139 diff2_2_or2v0x05_0_b 0 2.9fF
C140 diff2_0_an2v0x05_0_vdd 0 110.2fF
C141 diff2_0_an2v0x05_0_vss 0 66.5fF

v_dd diff2_0_an2v0x05_0_vdd 0 5
v_ss diff2_0_an2v0x05_0_vss 0 0
v_c1 diff2_0_an2v0x05_0_b 0 DC 1 PULSE(0 5 1ns 0.1ns 0.1ns 30ns 60ns )
v_a1 diff2_0_xnr2v0x05_0_b 0 DC 1 PULSE(0 5 1ns 0.1ns 0.1ns 30ns 60ns )
v_b1 diff2_0_an2v0x05_1_b 0 DC 1 PULSE(0 5 1ns 0.1ns 0.1ns 30ns 60ns )
v_a2 diff2_1_xnr2v0x05_0_b 0 DC 1 PULSE(0 5 1ns 0.1ns 0.1ns 30ns 60ns )
v_b2 diff2_1_an2v0x05_1_b 0 DC 1 PULSE(0 5 1ns 0.1ns 0.1ns 30ns 60ns )
v_a3 diff2_2_xnr2v0x05_0_b 0 DC 1 PULSE(0 5 1ns 0.1ns 0.1ns 30ns 60ns )
v_b3 diff2_2_an2v0x05_1_b 0 DC 1 PULSE(0 5 1ns 0.1ns 0.1ns 30ns 60ns )

.tran 0.01ns 60ns

.control
run
setplot tran1
plot diff2_0_xor3v0x05_0_z diff2_1_xor3v0x05_0_z diff2_2_xor3v0x05_0_z diff2_2_or2v0x05_0_z
.endc

.end 
