* Tue Aug 30 09:29:45 CEST 2005
.subckt iv1v7x1 a vdd vss z 
*SPICE circuit <iv1v7x1> from XCircuit v3.20

m1 z a vss vss n w=9u l=2.3636u ad='9u*5u+12p' as='9u*5u+12p' pd='9u*2+14u' ps='9u*2+14u'
m2 z a vdd vdd p w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
.ends
