* Mon Aug 16 14:10:58 CEST 2004
.subckt iv1v0x8 a vdd vss z 
*SPICE circuit <iv1v0x8> from XCircuit v3.10

m1 z a vss vss n w=52u l=2.3636u ad='52u*5u+12p' as='52u*5u+12p' pd='52u*2+14u' ps='52u*2+14u'
m2 z a vdd vdd p w=104u l=2.3636u ad='104u*5u+12p' as='104u*5u+12p' pd='104u*2+14u' ps='104u*2+14u'
.ends
