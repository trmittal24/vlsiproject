* Tue Aug 10 11:21:08 CEST 2004
.subckt xaon22_x1 a1 a2 b1 b2 vdd vss z 
*SPICE circuit <xaon22_x1> from XCircuit v3.10

m1 bn b1 vdd vdd p w=35u l=2.3636u ad='35u*5u+12p' as='35u*5u+12p' pd='35u*2+14u' ps='35u*2+14u'
m2 an a2 vdd vdd p w=35u l=2.3636u ad='35u*5u+12p' as='35u*5u+12p' pd='35u*2+14u' ps='35u*2+14u'
m3 n3 b2 an vss n w=23u l=2.3636u ad='23u*5u+12p' as='23u*5u+12p' pd='23u*2+14u' ps='23u*2+14u'
m4 z b1 n3 vss n w=23u l=2.3636u ad='23u*5u+12p' as='23u*5u+12p' pd='23u*2+14u' ps='23u*2+14u'
m5 n4 b1 vss vss n w=23u l=2.3636u ad='23u*5u+12p' as='23u*5u+12p' pd='23u*2+14u' ps='23u*2+14u'
m6 bn b2 n4 vss n w=23u l=2.3636u ad='23u*5u+12p' as='23u*5u+12p' pd='23u*2+14u' ps='23u*2+14u'
m7 an a1 vdd vdd p w=35u l=2.3636u ad='35u*5u+12p' as='35u*5u+12p' pd='35u*2+14u' ps='35u*2+14u'
m8 n2 a1 vss vss n w=33u l=2.3636u ad='33u*5u+12p' as='33u*5u+12p' pd='33u*2+14u' ps='33u*2+14u'
m9 an a2 n2 vss n w=33u l=2.3636u ad='33u*5u+12p' as='33u*5u+12p' pd='33u*2+14u' ps='33u*2+14u'
m10 z bn n1 vss n w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m11 z bn an vdd p w=35u l=2.3636u ad='35u*5u+12p' as='35u*5u+12p' pd='35u*2+14u' ps='35u*2+14u'
m12 n1 an vss vss n w=18u l=2.3636u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m13 bn b2 vdd vdd p w=35u l=2.3636u ad='35u*5u+12p' as='35u*5u+12p' pd='35u*2+14u' ps='35u*2+14u'
m14 z an bn vdd p w=35u l=2.3636u ad='35u*5u+12p' as='35u*5u+12p' pd='35u*2+14u' ps='35u*2+14u'
.ends
