* Thu Sep  1 18:58:43 CEST 2005
.subckt nr2v1x1 a b vdd vss z 
*SPICE circuit <nr2v1x1> from XCircuit v3.10

m1 z a vss vss n w=14u l=2.3636u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m2 n1 a vdd vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m3 z b vss vss n w=14u l=2.3636u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m4 z b n1 vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
.ends
