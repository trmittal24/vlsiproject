* Wed Apr  5 08:58:32 CEST 2006
.subckt bf1v0x12 a vdd vss z 
*SPICE circuit <bf1v0x12> from XCircuit v3.20

m1 an a vss vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m2 an a vdd vdd p w=60u l=2u ad='60u*5u+12p' as='60u*5u+12p' pd='60u*2+14u' ps='60u*2+14u'
m3 z an vss vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m4 z an vdd vdd p w=160u l=2u ad='160u*5u+12p' as='160u*5u+12p' pd='160u*2+14u' ps='160u*2+14u'
.ends
