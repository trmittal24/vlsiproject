* Spice description of nr2v0x2
* Spice driver version 134999461
* Date 17/05/2007 at  9:25:43
* wsclib 0.13um values
.subckt nr2v0x2 a b vdd vss z
M01 01    a     vdd   vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M02 vdd   a     05    vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M03 z     a     vss   vss n  L=0.12U  W=0.825U AS=0.218625P AD=0.218625P PS=2.18U   PD=2.18U
M04 z     b     01    vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M05 05    b     z     vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M06 vss   b     z     vss n  L=0.12U  W=0.825U AS=0.218625P AD=0.218625P PS=2.18U   PD=2.18U
C3  a     vss   0.682f
C4  b     vss   0.462f
C1  z     vss   0.672f
.ends
