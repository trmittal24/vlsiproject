* Mon Aug 16 14:10:59 CEST 2004
.subckt nr2v0x2 a b vdd vss z 
*SPICE circuit <nr2v0x2> from XCircuit v3.10

m1 z a vss vss n w=15u l=2.3636u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m2 n1 a vdd vdd p w=54u l=2.3636u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
m3 z b vss vss n w=15u l=2.3636u ad='15u*5u+12p' as='15u*5u+12p' pd='15u*2+14u' ps='15u*2+14u'
m4 z b n1 vdd p w=54u l=2.3636u ad='54u*5u+12p' as='54u*5u+12p' pd='54u*2+14u' ps='54u*2+14u'
.ends
