* Spice description of nd2_x05
* Spice driver version 134999461
* Date 31/05/2007 at 21:34:20
* vxlib 0.13um values
.subckt nd2_x05 a b vdd vss z
M1  z     b     vdd   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M2  vdd   a     z     vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M3  z     b     n1    vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
M4  n1    a     vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
C4  a     vss   0.499f
C5  b     vss   0.502f
C2  z     vss   0.846f
.ends
