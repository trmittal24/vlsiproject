* Tue Aug 10 11:21:07 CEST 2004
.subckt cgi2_x1 a b c vdd vss z 
*SPICE circuit <cgi2_x1> from XCircuit v3.10

m1 n4 a vss vss n w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m2 z b n4 vss n w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m3 n3 b vss vss n w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m4 z c n3 vss n w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m5 z b n2 vdd p w=39u l=2u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m6 n2 a vdd vdd p w=39u l=2u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m7 z c n1 vdd p w=39u l=2u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m8 n1 b vdd vdd p w=39u l=2u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m9 n1 a vdd vdd p w=39u l=2u ad='39u*5u+12p' as='39u*5u+12p' pd='39u*2+14u' ps='39u*2+14u'
m10 n3 a vss vss n w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
.ends
