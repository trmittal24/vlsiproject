* Spice description of nd3abv0x05
* Spice driver version 134999461
* Date 17/05/2007 at  9:21:54
* wsclib 0.13um values
.subckt nd3abv0x05 a b c vdd vss z
M01 06    b     03    vdd p  L=0.12U  W=0.825U AS=0.218625P AD=0.218625P PS=2.18U   PD=2.18U
M02 vss   b     06    vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M03 03    a     vdd   vdd p  L=0.12U  W=0.825U AS=0.218625P AD=0.218625P PS=2.18U   PD=2.18U
M04 06    a     vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M05 vdd   06    z     vdd p  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M06 vss   06    n2    vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M07 z     c     vdd   vdd p  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M08 n2    c     z     vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
C5  06    vss   0.601f
C7  a     vss   0.534f
C6  b     vss   0.630f
C4  c     vss   0.419f
C1  z     vss   0.595f
.ends
