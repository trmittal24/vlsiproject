* Tue Feb 20 08:57:11 CET 2007
.subckt iv1v0x8 a vdd vss z
*SPICE circuit <iv1v0x8> from XCircuit v3.4 rev 26

m1 z a vss vss n w=72u l=2.3636u ad='72u*5u+12p' as='72u*5u+12p' pd='72u*2+14u' ps='72u*2+14u'
m2 z a vdd vdd p w=104u l=2.3636u ad='104u*5u+12p' as='104u*5u+12p' pd='104u*2+14u' ps='104u*2+14u'
.ends
