* Spice description of buf_x4
* Spice driver version 134999461
* Date 21/07/2007 at 19:29:06
* sxlib 0.13um values
.subckt buf_x4 i q vdd vss
Mtr_00001 sig3  i     vss   vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00002 vss   sig3  q     vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00003 q     sig3  vss   vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00004 vdd   i     sig3  vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00005 vdd   sig3  q     vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00006 q     sig3  vdd   vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
C5  i     vss   0.981f
C2  q     vss   0.871f
C3  sig3  vss   0.789f
.ends
