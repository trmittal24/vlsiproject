* Tue Aug 10 11:21:07 CEST 2004
.subckt oai21_x2 a1 a2 b vdd vss z 
*SPICE circuit <oai21_x2> from XCircuit v3.10

m1 n1 a1 vdd vdd p w=76u l=2.3636u ad='76u*5u+12p' as='76u*5u+12p' pd='76u*2+14u' ps='76u*2+14u'
m2 z b vdd vdd p w=38u l=2.3636u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m3 n2 a2 vss vss n w=32u l=2.3636u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m4 n2 a1 vss vss n w=32u l=2.3636u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m5 z b n2 vss n w=32u l=2.3636u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m6 z a2 n1 vdd p w=76u l=2.3636u ad='76u*5u+12p' as='76u*5u+12p' pd='76u*2+14u' ps='76u*2+14u'
.ends
