* Spice description of aoi22v0x1
* Spice driver version 134999461
* Date 17/05/2007 at  9:01:32
* vsclib 0.13um values
.subckt aoi22v0x1 a1 a2 b1 b2 vdd vss z
M01 n3    a1    vdd   vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M02 vss   a1    sig6  vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M03 vdd   a2    n3    vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M04 sig6  a2    z     vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M05 z     b1    n3    vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M06 sig3  b1    vss   vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M07 n3    b2    z     vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M08 z     b2    sig3  vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
C7  a1    vss   0.525f
C8  a2    vss   0.477f
C4  b1    vss   0.417f
C5  b2    vss   0.422f
C9  n3    vss   0.305f
C2  z     vss   0.750f
.ends
