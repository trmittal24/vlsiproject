magic
tech scmos
timestamp 1520746549
<< pwell >>
rect -153 -31 295 5
<< nwell >>
rect -153 5 295 49
<< polysilicon >>
rect -140 39 -138 43
rect -94 41 -38 43
rect -94 33 -92 41
rect -84 33 -82 37
rect -74 33 -72 37
rect -67 33 -65 41
rect -57 33 -55 37
rect -50 33 -48 37
rect -130 25 -128 30
rect -111 27 -109 32
rect -104 27 -102 32
rect -140 7 -138 11
rect -130 8 -128 11
rect -130 7 -115 8
rect -140 6 -134 7
rect -130 6 -120 7
rect -140 2 -139 6
rect -135 2 -134 6
rect -140 1 -134 2
rect -122 3 -120 6
rect -116 3 -115 7
rect -122 2 -115 3
rect -140 -3 -138 1
rect -122 -1 -120 2
rect -111 -8 -109 21
rect -104 17 -102 21
rect -104 16 -98 17
rect -104 12 -103 16
rect -99 12 -98 16
rect -104 11 -98 12
rect -94 7 -92 21
rect -104 5 -92 7
rect -104 -8 -102 5
rect -84 2 -82 21
rect -74 17 -72 27
rect -78 16 -72 17
rect -78 12 -77 16
rect -73 12 -72 16
rect -78 11 -72 12
rect -84 1 -78 2
rect -98 0 -92 1
rect -98 -4 -97 0
rect -93 -4 -92 0
rect -98 -5 -92 -4
rect -94 -8 -92 -5
rect -84 -3 -83 1
rect -79 -3 -78 1
rect -84 -4 -78 -3
rect -84 -8 -82 -4
rect -74 -8 -72 11
rect -67 7 -65 27
rect -40 31 -38 41
rect 23 39 25 43
rect 33 39 35 43
rect 48 39 50 43
rect 58 39 60 43
rect -20 32 -18 37
rect -57 17 -55 20
rect -61 16 -55 17
rect -61 12 -60 16
rect -56 12 -55 16
rect -61 11 -55 12
rect -50 8 -48 20
rect -40 17 -38 20
rect -20 18 -18 22
rect -27 17 -18 18
rect -40 15 -32 17
rect -34 8 -32 15
rect -27 13 -26 17
rect -22 13 -18 17
rect -27 12 -18 13
rect -50 7 -44 8
rect -67 5 -55 7
rect -67 0 -61 1
rect -67 -4 -66 0
rect -62 -4 -61 0
rect -67 -5 -61 -4
rect -67 -8 -65 -5
rect -57 -8 -55 5
rect -50 3 -49 7
rect -45 3 -44 7
rect -50 2 -44 3
rect -34 7 -28 8
rect -34 3 -33 7
rect -29 3 -28 7
rect -34 2 -28 3
rect -50 -8 -48 2
rect -30 -1 -28 2
rect -20 -1 -18 12
rect 88 39 90 43
rect 98 39 100 43
rect 108 39 110 43
rect 118 39 120 43
rect 128 39 130 43
rect 156 39 158 43
rect 74 32 80 33
rect 68 24 70 29
rect 74 28 75 32
rect 79 28 80 32
rect 74 27 80 28
rect 78 24 80 27
rect 202 41 258 43
rect 202 33 204 41
rect 212 33 214 37
rect 222 33 224 37
rect 229 33 231 41
rect 239 33 241 37
rect 246 33 248 37
rect 166 25 168 30
rect 185 27 187 32
rect 192 27 194 32
rect 23 8 25 11
rect 33 8 35 11
rect 48 8 50 11
rect 58 8 60 11
rect 12 7 54 8
rect 12 3 13 7
rect 17 6 54 7
rect 17 3 24 6
rect 12 2 24 3
rect 12 -1 14 2
rect 22 -1 24 2
rect 42 -1 44 6
rect 52 -1 54 6
rect 58 7 64 8
rect 58 3 59 7
rect 63 3 64 7
rect 68 6 70 11
rect 78 6 80 11
rect 88 8 90 11
rect 98 8 100 11
rect 108 8 110 11
rect 88 7 100 8
rect 68 4 83 6
rect 58 2 64 3
rect 62 -1 64 2
rect 69 -1 71 4
rect 81 -1 83 4
rect 88 3 89 7
rect 93 6 100 7
rect 104 7 110 8
rect 93 3 94 6
rect 88 2 94 3
rect 104 3 105 7
rect 109 3 110 7
rect 104 2 110 3
rect 118 8 120 11
rect 128 8 130 11
rect 118 7 130 8
rect 118 3 125 7
rect 129 3 130 7
rect 118 2 130 3
rect 88 -1 90 2
rect 118 -1 120 2
rect 128 -1 130 2
rect 156 7 158 11
rect 166 8 168 11
rect 166 7 181 8
rect 156 6 162 7
rect 166 6 176 7
rect 156 2 157 6
rect 161 2 162 6
rect 156 1 162 2
rect 174 3 176 6
rect 180 3 181 7
rect 174 2 181 3
rect -122 -13 -120 -8
rect -30 -12 -28 -7
rect -20 -13 -18 -8
rect -140 -20 -138 -17
rect -111 -20 -109 -14
rect -104 -19 -102 -14
rect -140 -22 -109 -20
rect -94 -23 -92 -14
rect -84 -19 -82 -14
rect -74 -19 -72 -14
rect -67 -23 -65 -14
rect -57 -19 -55 -14
rect -50 -19 -48 -14
rect 12 -16 14 -12
rect -94 -25 -65 -23
rect 22 -23 24 -18
rect 42 -20 44 -15
rect 52 -20 54 -15
rect 62 -25 64 -20
rect 69 -25 71 -20
rect 156 -3 158 1
rect 174 -1 176 2
rect 118 -19 120 -15
rect 128 -19 130 -15
rect 185 -8 187 21
rect 192 17 194 21
rect 192 16 198 17
rect 192 12 193 16
rect 197 12 198 16
rect 192 11 198 12
rect 202 7 204 21
rect 192 5 204 7
rect 192 -8 194 5
rect 212 2 214 21
rect 222 17 224 27
rect 218 16 224 17
rect 218 12 219 16
rect 223 12 224 16
rect 218 11 224 12
rect 212 1 218 2
rect 198 0 204 1
rect 198 -4 199 0
rect 203 -4 204 0
rect 198 -5 204 -4
rect 202 -8 204 -5
rect 212 -3 213 1
rect 217 -3 218 1
rect 212 -4 218 -3
rect 212 -8 214 -4
rect 222 -8 224 11
rect 229 7 231 27
rect 256 31 258 41
rect 276 32 278 37
rect 239 17 241 20
rect 235 16 241 17
rect 235 12 236 16
rect 240 12 241 16
rect 235 11 241 12
rect 246 8 248 20
rect 256 17 258 20
rect 276 18 278 22
rect 269 17 278 18
rect 256 15 264 17
rect 262 8 264 15
rect 269 13 270 17
rect 274 13 278 17
rect 269 12 278 13
rect 246 7 252 8
rect 229 5 241 7
rect 229 0 235 1
rect 229 -4 230 0
rect 234 -4 235 0
rect 229 -5 235 -4
rect 229 -8 231 -5
rect 239 -8 241 5
rect 246 3 247 7
rect 251 3 252 7
rect 246 2 252 3
rect 262 7 268 8
rect 262 3 263 7
rect 267 3 268 7
rect 262 2 268 3
rect 246 -8 248 2
rect 266 -1 268 2
rect 276 -1 278 12
rect 174 -13 176 -8
rect 266 -12 268 -7
rect 276 -13 278 -8
rect 81 -25 83 -20
rect 88 -25 90 -20
rect 156 -20 158 -17
rect 185 -20 187 -14
rect 192 -19 194 -14
rect 156 -22 187 -20
rect 202 -23 204 -14
rect 212 -19 214 -14
rect 222 -19 224 -14
rect 229 -23 231 -14
rect 239 -19 241 -14
rect 246 -19 248 -14
rect 202 -25 231 -23
<< ndiffusion >>
rect -129 -2 -122 -1
rect -147 -4 -140 -3
rect -147 -8 -146 -4
rect -142 -8 -140 -4
rect -147 -9 -140 -8
rect -145 -17 -140 -9
rect -138 -11 -133 -3
rect -129 -6 -128 -2
rect -124 -6 -122 -2
rect -129 -7 -122 -6
rect -127 -8 -122 -7
rect -120 -8 -113 -1
rect -37 -2 -30 -1
rect -37 -6 -36 -2
rect -32 -6 -30 -2
rect -37 -7 -30 -6
rect -28 -2 -20 -1
rect -28 -6 -26 -2
rect -22 -6 -20 -2
rect -28 -7 -20 -6
rect -138 -12 -131 -11
rect -138 -16 -136 -12
rect -132 -16 -131 -12
rect -118 -9 -111 -8
rect -118 -13 -117 -9
rect -113 -13 -111 -9
rect -118 -14 -111 -13
rect -109 -14 -104 -8
rect -102 -9 -94 -8
rect -102 -13 -100 -9
rect -96 -13 -94 -9
rect -102 -14 -94 -13
rect -92 -9 -84 -8
rect -92 -13 -90 -9
rect -86 -13 -84 -9
rect -92 -14 -84 -13
rect -82 -9 -74 -8
rect -82 -13 -80 -9
rect -76 -13 -74 -9
rect -82 -14 -74 -13
rect -72 -14 -67 -8
rect -65 -9 -57 -8
rect -65 -13 -63 -9
rect -59 -13 -57 -9
rect -65 -14 -57 -13
rect -55 -14 -50 -8
rect -48 -9 -41 -8
rect -48 -13 -46 -9
rect -42 -13 -41 -9
rect -26 -8 -20 -7
rect -18 -2 -11 -1
rect -18 -6 -16 -2
rect -12 -6 -11 -2
rect -18 -8 -11 -6
rect 5 -7 12 -1
rect 5 -11 6 -7
rect 10 -11 12 -7
rect 5 -12 12 -11
rect 14 -2 22 -1
rect 14 -6 16 -2
rect 20 -6 22 -2
rect 14 -12 22 -6
rect -48 -14 -41 -13
rect -138 -17 -131 -16
rect 17 -18 22 -12
rect 24 -13 31 -1
rect 24 -17 26 -13
rect 30 -17 31 -13
rect 35 -2 42 -1
rect 35 -6 36 -2
rect 40 -6 42 -2
rect 35 -9 42 -6
rect 35 -13 36 -9
rect 40 -13 42 -9
rect 35 -15 42 -13
rect 44 -2 52 -1
rect 44 -6 46 -2
rect 50 -6 52 -2
rect 44 -15 52 -6
rect 54 -2 62 -1
rect 54 -6 56 -2
rect 60 -6 62 -2
rect 54 -9 62 -6
rect 54 -13 56 -9
rect 60 -13 62 -9
rect 54 -15 62 -13
rect 24 -18 31 -17
rect 57 -20 62 -15
rect 64 -20 69 -1
rect 71 -19 81 -1
rect 71 -20 74 -19
rect 73 -23 74 -20
rect 78 -20 81 -19
rect 83 -20 88 -1
rect 90 -8 95 -1
rect 90 -9 97 -8
rect 90 -13 92 -9
rect 96 -13 97 -9
rect 90 -14 97 -13
rect 90 -20 95 -14
rect 111 -10 118 -1
rect 111 -14 112 -10
rect 116 -14 118 -10
rect 111 -15 118 -14
rect 120 -2 128 -1
rect 120 -6 122 -2
rect 126 -6 128 -2
rect 120 -9 128 -6
rect 120 -13 122 -9
rect 126 -13 128 -9
rect 120 -15 128 -13
rect 130 -10 137 -1
rect 167 -2 174 -1
rect 149 -4 156 -3
rect 149 -8 150 -4
rect 154 -8 156 -4
rect 149 -9 156 -8
rect 130 -14 132 -10
rect 136 -14 137 -10
rect 130 -15 137 -14
rect 151 -17 156 -9
rect 158 -11 163 -3
rect 167 -6 168 -2
rect 172 -6 174 -2
rect 167 -7 174 -6
rect 169 -8 174 -7
rect 176 -8 183 -1
rect 259 -2 266 -1
rect 259 -6 260 -2
rect 264 -6 266 -2
rect 259 -7 266 -6
rect 268 -2 276 -1
rect 268 -6 270 -2
rect 274 -6 276 -2
rect 268 -7 276 -6
rect 158 -12 165 -11
rect 158 -16 160 -12
rect 164 -16 165 -12
rect 178 -9 185 -8
rect 178 -13 179 -9
rect 183 -13 185 -9
rect 178 -14 185 -13
rect 187 -14 192 -8
rect 194 -9 202 -8
rect 194 -13 196 -9
rect 200 -13 202 -9
rect 194 -14 202 -13
rect 204 -9 212 -8
rect 204 -13 206 -9
rect 210 -13 212 -9
rect 204 -14 212 -13
rect 214 -9 222 -8
rect 214 -13 216 -9
rect 220 -13 222 -9
rect 214 -14 222 -13
rect 224 -14 229 -8
rect 231 -9 239 -8
rect 231 -13 233 -9
rect 237 -13 239 -9
rect 231 -14 239 -13
rect 241 -14 246 -8
rect 248 -9 255 -8
rect 248 -13 250 -9
rect 254 -13 255 -9
rect 270 -8 276 -7
rect 278 -2 285 -1
rect 278 -6 280 -2
rect 284 -6 285 -2
rect 278 -8 285 -6
rect 248 -14 255 -13
rect 158 -17 165 -16
rect 78 -23 79 -20
rect 73 -24 79 -23
<< pdiffusion >>
rect -145 25 -140 39
rect -147 23 -140 25
rect -147 19 -146 23
rect -142 19 -140 23
rect -147 16 -140 19
rect -147 12 -146 16
rect -142 12 -140 16
rect -147 11 -140 12
rect -138 38 -131 39
rect -138 34 -136 38
rect -132 34 -131 38
rect -138 33 -131 34
rect -138 25 -132 33
rect -99 27 -94 33
rect -119 26 -111 27
rect -138 24 -130 25
rect -138 20 -136 24
rect -132 20 -130 24
rect -138 11 -130 20
rect -128 17 -123 25
rect -119 22 -118 26
rect -114 22 -111 26
rect -119 21 -111 22
rect -109 21 -104 27
rect -102 26 -94 27
rect -102 22 -100 26
rect -96 22 -94 26
rect -102 21 -94 22
rect -92 26 -84 33
rect -92 22 -90 26
rect -86 22 -84 26
rect -92 21 -84 22
rect -82 32 -74 33
rect -82 28 -80 32
rect -76 28 -74 32
rect -82 27 -74 28
rect -72 27 -67 33
rect -65 32 -57 33
rect -65 28 -63 32
rect -59 28 -57 32
rect -65 27 -57 28
rect -82 21 -76 27
rect -128 16 -121 17
rect -128 12 -126 16
rect -122 12 -121 16
rect -128 11 -121 12
rect -62 20 -57 27
rect -55 20 -50 33
rect -48 31 -43 33
rect -27 31 -20 32
rect -48 30 -40 31
rect -48 26 -46 30
rect -42 26 -40 30
rect -48 20 -40 26
rect -38 26 -33 31
rect -27 27 -26 31
rect -22 27 -20 31
rect -38 25 -31 26
rect -38 21 -36 25
rect -32 21 -31 25
rect -27 22 -20 27
rect -18 28 -13 32
rect -18 27 -11 28
rect -18 23 -16 27
rect -12 23 -11 27
rect -18 22 -11 23
rect -38 20 -31 21
rect 16 38 23 39
rect 16 34 17 38
rect 21 34 23 38
rect 16 31 23 34
rect 16 27 17 31
rect 21 27 23 31
rect 16 11 23 27
rect 25 23 33 39
rect 25 19 27 23
rect 31 19 33 23
rect 25 16 33 19
rect 25 12 27 16
rect 31 12 33 16
rect 25 11 33 12
rect 35 38 48 39
rect 35 34 39 38
rect 43 34 48 38
rect 35 31 48 34
rect 35 27 39 31
rect 43 27 48 31
rect 35 11 48 27
rect 50 31 58 39
rect 50 27 52 31
rect 56 27 58 31
rect 50 24 58 27
rect 50 20 52 24
rect 56 20 58 24
rect 50 11 58 20
rect 60 24 65 39
rect 83 24 88 39
rect 60 23 68 24
rect 60 19 62 23
rect 66 19 68 23
rect 60 16 68 19
rect 60 12 62 16
rect 66 12 68 16
rect 60 11 68 12
rect 70 16 78 24
rect 70 12 72 16
rect 76 12 78 16
rect 70 11 78 12
rect 80 23 88 24
rect 80 19 82 23
rect 86 19 88 23
rect 80 11 88 19
rect 90 32 98 39
rect 90 28 92 32
rect 96 28 98 32
rect 90 16 98 28
rect 90 12 92 16
rect 96 12 98 16
rect 90 11 98 12
rect 100 31 108 39
rect 100 27 102 31
rect 106 27 108 31
rect 100 24 108 27
rect 100 20 102 24
rect 106 20 108 24
rect 100 11 108 20
rect 110 23 118 39
rect 110 19 112 23
rect 116 19 118 23
rect 110 16 118 19
rect 110 12 112 16
rect 116 12 118 16
rect 110 11 118 12
rect 120 38 128 39
rect 120 34 122 38
rect 126 34 128 38
rect 120 31 128 34
rect 120 27 122 31
rect 126 27 128 31
rect 120 11 128 27
rect 130 24 135 39
rect 151 25 156 39
rect 130 23 137 24
rect 130 19 132 23
rect 136 19 137 23
rect 130 16 137 19
rect 130 12 132 16
rect 136 12 137 16
rect 130 11 137 12
rect 149 23 156 25
rect 149 19 150 23
rect 154 19 156 23
rect 149 16 156 19
rect 149 12 150 16
rect 154 12 156 16
rect 149 11 156 12
rect 158 38 165 39
rect 158 34 160 38
rect 164 34 165 38
rect 158 33 165 34
rect 158 25 164 33
rect 197 27 202 33
rect 177 26 185 27
rect 158 24 166 25
rect 158 20 160 24
rect 164 20 166 24
rect 158 11 166 20
rect 168 17 173 25
rect 177 22 178 26
rect 182 22 185 26
rect 177 21 185 22
rect 187 21 192 27
rect 194 26 202 27
rect 194 22 196 26
rect 200 22 202 26
rect 194 21 202 22
rect 204 26 212 33
rect 204 22 206 26
rect 210 22 212 26
rect 204 21 212 22
rect 214 32 222 33
rect 214 28 216 32
rect 220 28 222 32
rect 214 27 222 28
rect 224 27 229 33
rect 231 32 239 33
rect 231 28 233 32
rect 237 28 239 32
rect 231 27 239 28
rect 214 21 220 27
rect 168 16 175 17
rect 168 12 170 16
rect 174 12 175 16
rect 168 11 175 12
rect 234 20 239 27
rect 241 20 246 33
rect 248 31 253 33
rect 269 31 276 32
rect 248 30 256 31
rect 248 26 250 30
rect 254 26 256 30
rect 248 20 256 26
rect 258 26 263 31
rect 269 27 270 31
rect 274 27 276 31
rect 258 25 265 26
rect 258 21 260 25
rect 264 21 265 25
rect 269 22 276 27
rect 278 28 283 32
rect 278 27 285 28
rect 278 23 280 27
rect 284 23 285 27
rect 278 22 285 23
rect 258 20 265 21
<< metal1 >>
rect -151 41 293 45
rect -151 38 -122 41
rect -151 37 -136 38
rect -132 37 -122 38
rect -118 37 -112 41
rect -108 37 -31 41
rect -27 37 7 41
rect 11 38 72 41
rect 11 37 17 38
rect -136 24 -132 34
rect -147 23 -142 24
rect -147 19 -146 23
rect -118 26 -114 37
rect -80 32 -76 37
rect -80 27 -76 28
rect -68 28 -63 32
rect -59 28 -58 32
rect -47 30 -41 37
rect -90 26 -86 27
rect -118 21 -114 22
rect -111 22 -100 26
rect -96 22 -95 26
rect -136 19 -132 20
rect -147 16 -142 19
rect -147 12 -146 16
rect -142 12 -134 15
rect -147 11 -134 12
rect -128 12 -126 16
rect -122 12 -121 16
rect -147 -3 -143 11
rect -128 6 -124 12
rect -111 7 -107 22
rect -90 16 -86 22
rect -104 12 -103 16
rect -140 2 -139 6
rect -135 4 -124 6
rect -135 2 -128 4
rect -121 3 -120 7
rect -116 3 -105 7
rect -128 -2 -124 0
rect -147 -4 -142 -3
rect -147 -8 -146 -4
rect -128 -7 -124 -6
rect -147 -9 -142 -8
rect -117 -9 -113 -8
rect -136 -12 -132 -11
rect -136 -19 -132 -16
rect -109 -9 -105 3
rect -99 1 -95 16
rect -90 12 -77 16
rect -73 12 -72 16
rect -99 0 -93 1
rect -99 -4 -97 0
rect -99 -5 -93 -4
rect -90 -9 -86 12
rect -68 9 -64 28
rect -47 26 -46 30
rect -42 26 -41 30
rect -27 31 -21 37
rect -27 27 -26 31
rect -22 27 -21 31
rect 21 37 39 38
rect 17 31 21 34
rect -16 27 -12 28
rect -36 25 -32 26
rect -73 5 -64 9
rect -60 21 -36 23
rect 38 34 39 37
rect 43 37 72 38
rect 76 38 174 41
rect 76 37 122 38
rect 43 34 44 37
rect 38 31 44 34
rect 126 37 160 38
rect 38 27 39 31
rect 43 27 44 31
rect 52 31 75 32
rect 56 28 75 31
rect 79 28 92 32
rect 96 28 97 32
rect 101 31 106 32
rect 17 26 21 27
rect 52 24 56 27
rect -60 19 -32 21
rect -60 16 -56 19
rect -28 17 -22 23
rect -28 15 -26 17
rect -73 2 -69 5
rect -83 1 -69 2
rect -60 1 -56 12
rect -52 7 -46 15
rect -36 13 -26 15
rect -36 11 -22 13
rect -16 7 -12 23
rect 26 19 27 23
rect 31 20 52 23
rect 101 27 102 31
rect 101 24 106 27
rect 122 31 126 34
rect 122 26 126 27
rect 164 37 174 38
rect 178 37 184 41
rect 188 37 265 41
rect 269 37 293 41
rect 160 24 164 34
rect 101 23 102 24
rect 31 19 56 20
rect 61 19 62 23
rect 66 19 82 23
rect 86 20 102 23
rect 86 19 106 20
rect 111 23 116 24
rect 111 19 112 23
rect 26 16 31 19
rect -52 3 -49 7
rect -45 3 -42 7
rect -34 3 -33 7
rect -29 3 -16 7
rect -79 -3 -69 1
rect -83 -4 -69 -3
rect -109 -13 -100 -9
rect -96 -13 -95 -9
rect -117 -19 -113 -13
rect -90 -14 -86 -13
rect -80 -9 -76 -8
rect -73 -9 -69 -4
rect -66 0 -56 1
rect -62 -1 -56 0
rect -62 -2 -31 -1
rect -62 -4 -36 -2
rect -66 -5 -36 -4
rect -37 -6 -36 -5
rect -32 -6 -31 -2
rect -26 -2 -22 -1
rect -73 -13 -63 -9
rect -59 -13 -58 -9
rect -47 -13 -46 -9
rect -42 -13 -41 -9
rect -80 -19 -76 -13
rect -47 -19 -41 -13
rect -26 -19 -22 -6
rect -16 -2 -12 3
rect 5 8 9 16
rect 26 12 27 16
rect 61 16 66 19
rect 111 16 116 19
rect 132 23 137 24
rect 136 19 137 23
rect 132 16 137 19
rect 61 15 62 16
rect 26 11 31 12
rect 37 12 62 15
rect 37 11 66 12
rect 71 12 72 16
rect 76 12 77 16
rect 5 7 17 8
rect 5 3 13 7
rect 5 2 17 3
rect 26 -2 30 11
rect 37 4 41 11
rect 71 7 77 12
rect 91 12 92 16
rect 96 15 97 16
rect 96 12 106 15
rect 111 12 112 16
rect 116 12 132 16
rect 136 12 137 16
rect 149 23 154 24
rect 149 19 150 23
rect 178 26 182 37
rect 216 32 220 37
rect 216 27 220 28
rect 228 28 233 32
rect 237 28 238 32
rect 249 30 255 37
rect 206 26 210 27
rect 178 21 182 22
rect 185 22 196 26
rect 200 22 201 26
rect 160 19 164 20
rect 149 16 154 19
rect 149 12 150 16
rect 154 12 162 15
rect 91 11 106 12
rect 102 7 106 11
rect 37 -2 41 0
rect 15 -6 16 -2
rect 20 -6 30 -2
rect 35 -6 36 -2
rect 40 -6 41 -2
rect 45 3 59 7
rect 63 3 89 7
rect 93 3 96 7
rect 102 3 105 7
rect 109 3 110 7
rect 45 -2 51 3
rect 92 -1 96 3
rect 115 -1 119 12
rect 149 11 162 12
rect 168 12 170 16
rect 174 12 175 16
rect 124 7 137 8
rect 124 3 125 7
rect 129 3 137 7
rect 149 3 153 11
rect 168 6 172 12
rect 185 7 189 22
rect 206 16 210 22
rect 192 12 193 16
rect 133 0 153 3
rect 156 2 157 6
rect 161 4 172 6
rect 161 2 168 4
rect 45 -6 46 -2
rect 50 -6 51 -2
rect 56 -2 60 -1
rect 92 -2 126 -1
rect 92 -5 122 -2
rect -16 -7 -12 -6
rect 6 -7 10 -6
rect 6 -19 10 -11
rect 35 -9 41 -6
rect 56 -9 60 -6
rect 133 -6 137 0
rect 149 -3 153 0
rect 175 3 176 7
rect 180 3 191 7
rect 168 -2 172 0
rect 149 -4 154 -3
rect 122 -9 126 -6
rect 149 -8 150 -4
rect 168 -7 172 -6
rect 149 -9 154 -8
rect 179 -9 183 -8
rect 26 -13 30 -12
rect 35 -13 36 -9
rect 40 -13 56 -9
rect 60 -13 92 -9
rect 96 -13 98 -9
rect 112 -10 116 -9
rect 26 -19 30 -17
rect 122 -14 126 -13
rect 131 -14 132 -10
rect 136 -14 137 -10
rect 112 -19 116 -14
rect 131 -19 137 -14
rect 160 -12 164 -11
rect 160 -19 164 -16
rect 187 -9 191 3
rect 197 1 201 16
rect 206 12 219 16
rect 223 12 224 16
rect 197 0 203 1
rect 197 -4 199 0
rect 197 -5 203 -4
rect 206 -9 210 12
rect 228 9 232 28
rect 249 26 250 30
rect 254 26 255 30
rect 269 31 275 37
rect 269 27 270 31
rect 274 27 275 31
rect 280 27 284 28
rect 260 25 264 26
rect 223 5 232 9
rect 236 21 260 23
rect 236 19 264 21
rect 236 16 240 19
rect 268 17 274 23
rect 268 15 270 17
rect 223 2 227 5
rect 213 1 227 2
rect 236 1 240 12
rect 244 7 250 15
rect 260 13 270 15
rect 260 11 274 13
rect 280 7 284 23
rect 244 3 247 7
rect 251 3 254 7
rect 262 3 263 7
rect 267 3 284 7
rect 217 -3 227 1
rect 213 -4 227 -3
rect 187 -13 196 -9
rect 200 -13 201 -9
rect 179 -19 183 -13
rect 206 -14 210 -13
rect 216 -9 220 -8
rect 223 -9 227 -4
rect 230 0 240 1
rect 234 -1 240 0
rect 234 -2 265 -1
rect 234 -4 260 -2
rect 230 -5 260 -4
rect 259 -6 260 -5
rect 264 -6 265 -2
rect 270 -2 274 -1
rect 223 -13 233 -9
rect 237 -13 238 -9
rect 249 -13 250 -9
rect 254 -13 255 -9
rect 216 -19 220 -13
rect 249 -19 255 -13
rect 270 -19 274 -6
rect 280 -2 284 3
rect 280 -7 284 -6
rect -151 -23 -30 -19
rect -26 -23 -19 -19
rect -15 -23 7 -19
rect 11 -23 74 -19
rect 78 -23 102 -19
rect 106 -23 266 -19
rect 270 -23 277 -19
rect 281 -23 293 -19
rect -151 -27 293 -23
<< metal2 >>
rect -42 0 -38 3
rect -12 3 37 4
rect -16 0 37 3
rect 254 0 258 3
rect -128 -3 -38 0
rect 168 -3 258 0
<< ntransistor >>
rect -140 -17 -138 -3
rect -122 -8 -120 -1
rect -30 -7 -28 -1
rect -111 -14 -109 -8
rect -104 -14 -102 -8
rect -94 -14 -92 -8
rect -84 -14 -82 -8
rect -74 -14 -72 -8
rect -67 -14 -65 -8
rect -57 -14 -55 -8
rect -50 -14 -48 -8
rect -20 -8 -18 -1
rect 12 -12 14 -1
rect 22 -18 24 -1
rect 42 -15 44 -1
rect 52 -15 54 -1
rect 62 -20 64 -1
rect 69 -20 71 -1
rect 81 -20 83 -1
rect 88 -20 90 -1
rect 118 -15 120 -1
rect 128 -15 130 -1
rect 156 -17 158 -3
rect 174 -8 176 -1
rect 266 -7 268 -1
rect 185 -14 187 -8
rect 192 -14 194 -8
rect 202 -14 204 -8
rect 212 -14 214 -8
rect 222 -14 224 -8
rect 229 -14 231 -8
rect 239 -14 241 -8
rect 246 -14 248 -8
rect 276 -8 278 -1
<< ptransistor >>
rect -140 11 -138 39
rect -130 11 -128 25
rect -111 21 -109 27
rect -104 21 -102 27
rect -94 21 -92 33
rect -84 21 -82 33
rect -74 27 -72 33
rect -67 27 -65 33
rect -57 20 -55 33
rect -50 20 -48 33
rect -40 20 -38 31
rect -20 22 -18 32
rect 23 11 25 39
rect 33 11 35 39
rect 48 11 50 39
rect 58 11 60 39
rect 68 11 70 24
rect 78 11 80 24
rect 88 11 90 39
rect 98 11 100 39
rect 108 11 110 39
rect 118 11 120 39
rect 128 11 130 39
rect 156 11 158 39
rect 166 11 168 25
rect 185 21 187 27
rect 192 21 194 27
rect 202 21 204 33
rect 212 21 214 33
rect 222 27 224 33
rect 229 27 231 33
rect 239 20 241 33
rect 246 20 248 33
rect 256 20 258 31
rect 276 22 278 32
<< polycontact >>
rect -139 2 -135 6
rect -120 3 -116 7
rect -103 12 -99 16
rect -77 12 -73 16
rect -97 -4 -93 0
rect -83 -3 -79 1
rect -60 12 -56 16
rect -26 13 -22 17
rect -66 -4 -62 0
rect -49 3 -45 7
rect -33 3 -29 7
rect 75 28 79 32
rect 13 3 17 7
rect 59 3 63 7
rect 89 3 93 7
rect 105 3 109 7
rect 125 3 129 7
rect 157 2 161 6
rect 176 3 180 7
rect 193 12 197 16
rect 219 12 223 16
rect 199 -4 203 0
rect 213 -3 217 1
rect 236 12 240 16
rect 270 13 274 17
rect 230 -4 234 0
rect 247 3 251 7
rect 263 3 267 7
<< ndcontact >>
rect -146 -8 -142 -4
rect -128 -6 -124 -2
rect -36 -6 -32 -2
rect -26 -6 -22 -2
rect -136 -16 -132 -12
rect -117 -13 -113 -9
rect -100 -13 -96 -9
rect -90 -13 -86 -9
rect -80 -13 -76 -9
rect -63 -13 -59 -9
rect -46 -13 -42 -9
rect -16 -6 -12 -2
rect 6 -11 10 -7
rect 16 -6 20 -2
rect 26 -17 30 -13
rect 36 -6 40 -2
rect 36 -13 40 -9
rect 46 -6 50 -2
rect 56 -6 60 -2
rect 56 -13 60 -9
rect 74 -23 78 -19
rect 92 -13 96 -9
rect 112 -14 116 -10
rect 122 -6 126 -2
rect 122 -13 126 -9
rect 150 -8 154 -4
rect 132 -14 136 -10
rect 168 -6 172 -2
rect 260 -6 264 -2
rect 270 -6 274 -2
rect 160 -16 164 -12
rect 179 -13 183 -9
rect 196 -13 200 -9
rect 206 -13 210 -9
rect 216 -13 220 -9
rect 233 -13 237 -9
rect 250 -13 254 -9
rect 280 -6 284 -2
<< pdcontact >>
rect -146 19 -142 23
rect -146 12 -142 16
rect -136 34 -132 38
rect -136 20 -132 24
rect -118 22 -114 26
rect -100 22 -96 26
rect -90 22 -86 26
rect -80 28 -76 32
rect -63 28 -59 32
rect -126 12 -122 16
rect -46 26 -42 30
rect -26 27 -22 31
rect -36 21 -32 25
rect -16 23 -12 27
rect 17 34 21 38
rect 17 27 21 31
rect 27 19 31 23
rect 27 12 31 16
rect 39 34 43 38
rect 39 27 43 31
rect 52 27 56 31
rect 52 20 56 24
rect 62 19 66 23
rect 62 12 66 16
rect 72 12 76 16
rect 82 19 86 23
rect 92 28 96 32
rect 92 12 96 16
rect 102 27 106 31
rect 102 20 106 24
rect 112 19 116 23
rect 112 12 116 16
rect 122 34 126 38
rect 122 27 126 31
rect 132 19 136 23
rect 132 12 136 16
rect 150 19 154 23
rect 150 12 154 16
rect 160 34 164 38
rect 160 20 164 24
rect 178 22 182 26
rect 196 22 200 26
rect 206 22 210 26
rect 216 28 220 32
rect 233 28 237 32
rect 170 12 174 16
rect 250 26 254 30
rect 270 27 274 31
rect 260 21 264 25
rect 280 23 284 27
<< m2contact >>
rect -128 0 -124 4
rect -42 3 -38 7
rect -16 3 -12 7
rect 37 0 41 4
rect 168 0 172 4
rect 254 3 258 7
<< psubstratepcontact >>
rect -30 -23 -26 -19
rect -19 -23 -15 -19
rect 7 -23 11 -19
rect 102 -23 106 -19
rect 266 -23 270 -19
rect 277 -23 281 -19
<< nsubstratencontact >>
rect -122 37 -118 41
rect -112 37 -108 41
rect -31 37 -27 41
rect 7 37 11 41
rect 72 37 76 41
rect 174 37 178 41
rect 184 37 188 41
rect 265 37 269 41
<< psubstratepdiff >>
rect -37 -19 -8 -18
rect -37 -23 -30 -19
rect -26 -23 -19 -19
rect -15 -23 -8 -19
rect -37 -24 -8 -23
rect 6 -19 12 -18
rect 6 -23 7 -19
rect 11 -23 12 -19
rect 6 -24 12 -23
rect 101 -19 107 -3
rect 101 -23 102 -19
rect 106 -23 107 -19
rect 101 -24 107 -23
rect 259 -19 288 -18
rect 259 -23 266 -19
rect 270 -23 277 -19
rect 281 -23 288 -19
rect 259 -24 288 -23
<< nsubstratendiff >>
rect -127 41 -103 42
rect -127 37 -122 41
rect -118 37 -112 41
rect -108 37 -103 41
rect -127 36 -103 37
rect -32 41 -26 42
rect -32 37 -31 41
rect -27 37 -26 41
rect 6 41 12 42
rect 6 37 7 41
rect 11 37 12 41
rect 71 41 77 42
rect -32 36 -26 37
rect 6 13 12 37
rect 71 37 72 41
rect 76 37 77 41
rect 169 41 193 42
rect 71 36 77 37
rect 169 37 174 41
rect 178 37 184 41
rect 188 37 193 41
rect 169 36 193 37
rect 264 41 270 42
rect 264 37 265 41
rect 269 37 270 41
rect 264 36 270 37
<< labels >>
rlabel polycontact -137 4 -137 4 6 zn
rlabel polycontact -119 5 -119 5 6 n4
rlabel polycontact -95 -2 -95 -2 6 ci
rlabel polycontact -101 14 -101 14 6 ci
rlabel polycontact -81 -1 -81 -1 6 n1
rlabel polycontact -64 -2 -64 -2 6 ci
rlabel polycontact -58 14 -58 14 6 ci
rlabel polycontact -75 14 -75 14 6 n2
rlabel polycontact -31 5 -31 5 6 cn
rlabel metal1 -132 4 -132 4 6 zn
rlabel metal1 -126 4 -126 4 6 zn
rlabel metal1 -102 -11 -102 -11 6 n4
rlabel polycontact -96 -2 -96 -2 6 ci
rlabel metal1 -113 5 -113 5 6 n4
rlabel polycontact -100 14 -100 14 6 ci
rlabel metal1 -103 24 -103 24 6 n4
rlabel metal1 -77 -23 -77 -23 6 vss
rlabel metal1 -76 -1 -76 -1 6 n1
rlabel metal1 -81 14 -81 14 6 n2
rlabel metal1 -88 6 -88 6 6 n2
rlabel metal1 -77 41 -77 41 6 vdd
rlabel metal1 -66 -11 -66 -11 6 n1
rlabel m2contact -41 5 -41 5 6 d
rlabel metal1 -49 9 -49 9 6 d
rlabel metal1 -58 9 -58 9 6 ci
rlabel metal1 -63 30 -63 30 6 n1
rlabel metal1 -49 -3 -49 -3 6 ci
rlabel metal1 -23 5 -23 5 6 cn
rlabel metal1 -14 10 -14 10 6 cn
rlabel pdcontact -34 22 -34 22 6 ci
rlabel polycontact 91 5 91 5 6 an
rlabel polycontact 77 30 77 30 6 bn
rlabel polycontact 107 5 107 5 6 bn
rlabel metal1 47 -11 47 -11 6 z
rlabel metal1 22 -4 22 -4 6 bn
rlabel ndcontact 39 -3 39 -3 6 z
rlabel metal1 48 0 48 0 6 an
rlabel metal1 47 13 47 13 6 z
rlabel metal1 28 8 28 8 6 bn
rlabel metal1 54 25 54 25 6 bn
rlabel metal1 71 -23 71 -23 6 vss
rlabel metal1 79 -11 79 -11 6 z
rlabel metal1 71 -11 71 -11 6 z
rlabel metal1 63 -11 63 -11 6 z
rlabel metal1 55 -11 55 -11 6 z
rlabel metal1 55 13 55 13 6 z
rlabel pdcontact 63 13 63 13 6 z
rlabel metal1 74 9 74 9 6 an
rlabel metal1 79 21 79 21 6 z
rlabel metal1 71 21 71 21 6 z
rlabel metal1 71 41 71 41 6 vdd
rlabel ndcontact 95 -11 95 -11 6 z
rlabel metal1 87 -11 87 -11 6 z
rlabel metal1 104 9 104 9 6 bn
rlabel metal1 70 5 70 5 6 an
rlabel pdcontact 94 13 94 13 6 bn
rlabel metal1 87 21 87 21 6 z
rlabel metal1 103 25 103 25 6 z
rlabel metal1 95 21 95 21 6 z
rlabel metal1 74 30 74 30 6 bn
rlabel metal1 124 -8 124 -8 6 an
rlabel metal1 135 1 135 1 6 a
rlabel polycontact 127 5 127 5 6 a
rlabel metal1 134 18 134 18 6 an
rlabel metal1 124 14 124 14 6 an
rlabel metal1 113 18 113 18 6 an
rlabel polycontact 159 4 159 4 6 zn
rlabel polycontact 177 5 177 5 6 n4
rlabel polycontact 201 -2 201 -2 6 ci
rlabel polycontact 195 14 195 14 6 ci
rlabel polycontact 215 -1 215 -1 6 n1
rlabel polycontact 232 -2 232 -2 6 ci
rlabel polycontact 238 14 238 14 6 ci
rlabel polycontact 221 14 221 14 6 n2
rlabel polycontact 265 5 265 5 6 cn
rlabel metal1 164 4 164 4 6 zn
rlabel metal1 170 4 170 4 6 zn
rlabel metal1 194 -11 194 -11 6 n4
rlabel polycontact 200 -2 200 -2 6 ci
rlabel metal1 183 5 183 5 6 n4
rlabel polycontact 196 14 196 14 6 ci
rlabel metal1 193 24 193 24 6 n4
rlabel metal1 219 -23 219 -23 6 vss
rlabel metal1 220 -1 220 -1 6 n1
rlabel metal1 215 14 215 14 6 n2
rlabel metal1 208 6 208 6 6 n2
rlabel metal1 219 41 219 41 6 vdd
rlabel metal1 230 -11 230 -11 6 n1
rlabel m2contact 255 5 255 5 6 d
rlabel metal1 247 9 247 9 6 d
rlabel metal1 238 9 238 9 6 ci
rlabel metal1 233 30 233 30 6 n1
rlabel metal1 247 -3 247 -3 6 ci
rlabel metal1 273 5 273 5 6 cn
rlabel metal1 263 13 263 13 6 cp
rlabel metal1 271 17 271 17 6 cp
rlabel metal1 282 10 282 10 6 cn
rlabel pdcontact 262 22 262 22 6 ci
rlabel metal1 151 9 151 9 1 q0
rlabel metal1 159 13 159 13 1 q0
rlabel metal1 7 9 7 9 1 ud
rlabel polycontact 15 5 15 5 1 ud
rlabel metal1 -145 9 -145 9 1 q1
rlabel metal1 -137 13 -137 13 1 q1
rlabel metal1 -33 13 -33 13 1 cp1
rlabel polycontact -25 17 -25 17 1 cp1
<< end >>
