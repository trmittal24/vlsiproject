* Mon Sep 12 14:09:09 CEST 2005
.subckt or3v0x2 a b c vdd vss z 
*SPICE circuit <or3v0x2> from XCircuit v3.20

m1 zn c n2 vdd p w=42u l=2.3636u ad='42u*5u+12p' as='42u*5u+12p' pd='42u*2+14u' ps='42u*2+14u'
m2 n2 b n1 vdd p w=42u l=2.3636u ad='42u*5u+12p' as='42u*5u+12p' pd='42u*2+14u' ps='42u*2+14u'
m3 z zn vdd vdd p w=28u l=2.3636u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m4 z zn vss vss n w=14u l=2.3636u ad='14u*5u+12p' as='14u*5u+12p' pd='14u*2+14u' ps='14u*2+14u'
m5 zn a vss vss n w=8u l=2.3636u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
m6 zn b vss vss n w=8u l=2.3636u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
m7 zn c vss vss n w=8u l=2.3636u ad='8u*5u+12p' as='8u*5u+12p' pd='8u*2+14u' ps='8u*2+14u'
m8 n1 a vdd vdd p w=42u l=2.3636u ad='42u*5u+12p' as='42u*5u+12p' pd='42u*2+14u' ps='42u*2+14u'
.ends
