* Mon Aug 16 14:10:57 CEST 2004
.subckt an4v0x4 a b c d vdd vss z 
*SPICE circuit <an4v0x4> from XCircuit v3.10

m1 zn a vdd vdd p w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m2 zn b vdd vdd p w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m3 zn c vdd vdd p w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m4 zn d n3 vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m5 n3 c n2 vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m6 n2 b n1 vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
m7 z zn vss vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m8 z zn vdd vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m9 zn d vdd vdd p w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m10 n1 a vss vss n w=32u l=2u ad='32u*5u+12p' as='32u*5u+12p' pd='32u*2+14u' ps='32u*2+14u'
.ends
