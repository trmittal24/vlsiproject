* Tue Aug 10 11:21:07 CEST 2004
.subckt nr2_x2 a b vdd vss z 
*SPICE circuit <nr2_x2> from XCircuit v3.10

m1 z a vss vss n w=21u l=2.3636u ad='21u*5u+12p' as='21u*5u+12p' pd='21u*2+14u' ps='21u*2+14u'
m2 n1 a vdd vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
m3 z b vss vss n w=21u l=2.3636u ad='21u*5u+12p' as='21u*5u+12p' pd='21u*2+14u' ps='21u*2+14u'
m4 z b n1 vdd p w=78u l=2.3636u ad='78u*5u+12p' as='78u*5u+12p' pd='78u*2+14u' ps='78u*2+14u'
.ends
