* Tue Apr  4 18:58:30 CEST 2006
.subckt iv1v3x6 a vdd vss z 
*SPICE circuit <iv1v3x6> from XCircuit v3.20

m1 z a vss vss n w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
m2 z a vdd vdd p w=80u l=2u ad='80u*5u+12p' as='80u*5u+12p' pd='80u*2+14u' ps='80u*2+14u'
.ends
