* Mon Sep 12 14:09:07 CEST 2005
.subckt or3v0x05 a b c vdd vss z 
*SPICE circuit <or3v0x05> from XCircuit v3.20

m1 zn c n2 vdd p w=25u l=2.3636u ad='25u*5u+12p' as='25u*5u+12p' pd='25u*2+14u' ps='25u*2+14u'
m2 n2 b n1 vdd p w=25u l=2.3636u ad='25u*5u+12p' as='25u*5u+12p' pd='25u*2+14u' ps='25u*2+14u'
m3 z zn vdd vdd p w=12u l=2.3636u ad='12u*5u+12p' as='12u*5u+12p' pd='12u*2+14u' ps='12u*2+14u'
m4 z zn vss vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m5 zn a vss vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m6 zn b vss vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m7 zn c vss vss n w=6u l=2.3636u ad='6u*5u+12p' as='6u*5u+12p' pd='6u*2+14u' ps='6u*2+14u'
m8 n1 a vdd vdd p w=25u l=2.3636u ad='25u*5u+12p' as='25u*5u+12p' pd='25u*2+14u' ps='25u*2+14u'
.ends
