* Spice description of iv2_x2
* Spice driver version 134934782
* Date 15/09/2003 at 17:02:16
*
.subckt iv2_x2 a vdd vss z 
M1  vdd   a     z     vdd p  L=0.13U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U  
M2  vss   a     z     vss n  L=0.13U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U   
C4  a     vss   1.267f
C3  vdd   vss   0.847f
C2  z     vss   1.948f
.ends
