* Mon Aug 16 14:10:58 CEST 2004
.subckt iv1v1x4 a vdd vss z 
*SPICE circuit <iv1v1x4> from XCircuit v3.10

m1 z a vss vss n w=38u l=2.3636u ad='38u*5u+12p' as='38u*5u+12p' pd='38u*2+14u' ps='38u*2+14u'
m2 z a vdd vdd p w=56u l=2.3636u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
.ends
