* Spice description of vfeed7
* Spice driver version 134999461
* Date 22/07/2007 at 11:00:28
* vsxlib 0.13um values
.subckt vfeed7 vdd vss
.ends
