* Sat Aug 27 19:28:29 CEST 2005
.subckt nd2v5x4 a b vdd vss z 
*SPICE circuit <nd2v5x4> from XCircuit v3.20

m1 n1 a vss vss n w=36u l=2u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
m2 z a vdd vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
m3 z b n1 vss n w=36u l=2u ad='36u*5u+12p' as='36u*5u+12p' pd='36u*2+14u' ps='36u*2+14u'
m4 z b vdd vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
.ends
