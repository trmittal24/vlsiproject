* SPICE3 file created from totdiff2.ext - technology: scmos

.include t14y_tsmc_025_level3.txt
M1000 mux_0_vdd diff2_2_an2v0x2_2_zn diff2_2_an2v0x2_2_z mux_0_vdd pfet w=28u l=2u
+  ad=11922p pd=4362u as=166p ps=70u
M1001 diff2_2_an2v0x2_2_zn diff2_2_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1002 mux_0_vdd diff2_2_in_2c diff2_2_an2v0x2_2_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1003 mux_0_gnd diff2_2_an2v0x2_2_zn diff2_2_an2v0x2_2_z mux_0_gnd nfet w=14u l=2u
+  ad=8469p pd=3006u as=98p ps=42u
M1004 diff2_2_an2v0x2_2_a_24_13# diff2_2_an2v0x2_2_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1005 diff2_2_an2v0x2_2_zn diff2_2_in_2c diff2_2_an2v0x2_2_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1006 diff2_2_xor2v2x2_0_an diff2_2_xor2v2x2_0_bn mux_0_b2 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1007 mux_0_b2 diff2_2_xor2v2x2_0_bn diff2_2_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1008 diff2_2_xor2v2x2_0_bn diff2_2_xor2v2x2_0_an mux_0_b2 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1009 mux_0_b2 diff2_2_xor2v2x2_0_an diff2_2_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1010 diff2_2_xor2v2x2_0_bn diff2_2_in_2c mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1011 mux_0_vdd diff2_2_in_2c diff2_2_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1012 diff2_2_xor2v2x2_0_an diff2_2_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1013 mux_0_vdd diff2_2_an2v0x2_2_a diff2_2_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1014 diff2_2_xor2v2x2_0_a_13_13# diff2_2_xor2v2x2_0_an mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1015 mux_0_b2 diff2_2_xor2v2x2_0_bn diff2_2_xor2v2x2_0_a_13_13# mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1016 diff2_2_xor2v2x2_0_a_30_13# diff2_2_xor2v2x2_0_bn mux_0_b2 mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1017 mux_0_gnd diff2_2_xor2v2x2_0_an diff2_2_xor2v2x2_0_a_30_13# mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1018 diff2_2_xor2v2x2_0_bn diff2_2_in_2c mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1019 mux_0_b2 diff2_2_an2v0x2_2_a diff2_2_xor2v2x2_0_bn mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1020 diff2_2_xor2v2x2_0_an diff2_2_in_2c mux_0_b2 mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1021 mux_0_gnd diff2_2_an2v0x2_2_a diff2_2_xor2v2x2_0_an mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1022 mux_0_s diff2_2_or2v0x3_0_zn mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1023 mux_0_vdd diff2_2_or2v0x3_0_zn mux_0_s mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1024 diff2_2_or2v0x3_0_a_31_39# diff2_2_an2v0x2_1_z mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1025 diff2_2_or2v0x3_0_zn diff2_2_an2v0x2_0_z diff2_2_or2v0x3_0_a_31_39# mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1026 diff2_2_or2v0x3_0_a_48_39# diff2_2_an2v0x2_0_z diff2_2_or2v0x3_0_zn mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1027 mux_0_vdd diff2_2_an2v0x2_1_z diff2_2_or2v0x3_0_a_48_39# mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1028 mux_0_gnd diff2_2_or2v0x3_0_zn mux_0_s mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1029 diff2_2_or2v0x3_0_zn diff2_2_an2v0x2_1_z mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1030 mux_0_gnd diff2_2_an2v0x2_0_z diff2_2_or2v0x3_0_zn mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1031 mux_0_vdd diff2_2_an2v0x2_1_zn diff2_2_an2v0x2_1_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1032 diff2_2_an2v0x2_1_zn diff2_2_an2v0x2_1_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1033 mux_0_vdd diff2_2_in_b diff2_2_an2v0x2_1_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1034 mux_0_gnd diff2_2_an2v0x2_1_zn diff2_2_an2v0x2_1_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1035 diff2_2_an2v0x2_1_a_24_13# diff2_2_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1036 diff2_2_an2v0x2_1_zn diff2_2_in_b diff2_2_an2v0x2_1_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1037 mux_0_vdd diff2_2_an2v0x2_0_zn diff2_2_an2v0x2_0_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1038 diff2_2_an2v0x2_0_zn diff2_2_in_c mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1039 mux_0_vdd diff2_2_an2v0x2_0_b diff2_2_an2v0x2_0_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1040 mux_0_gnd diff2_2_an2v0x2_0_zn diff2_2_an2v0x2_0_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1041 diff2_2_an2v0x2_0_a_24_13# diff2_2_in_c mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1042 diff2_2_an2v0x2_0_zn diff2_2_an2v0x2_0_b diff2_2_an2v0x2_0_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1043 mux_0_vdd diff2_2_xnr2v8x05_0_zn diff2_2_an2v0x2_0_b mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1044 diff2_2_xnr2v8x05_0_an diff2_2_in_a mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1045 diff2_2_xnr2v8x05_0_zn diff2_2_xnr2v8x05_0_bn diff2_2_xnr2v8x05_0_an mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1046 diff2_2_xnr2v8x05_0_ai diff2_2_in_b diff2_2_xnr2v8x05_0_zn mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1047 mux_0_vdd diff2_2_xnr2v8x05_0_an diff2_2_xnr2v8x05_0_ai mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1048 diff2_2_xnr2v8x05_0_bn diff2_2_in_b mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1049 mux_0_gnd diff2_2_xnr2v8x05_0_zn diff2_2_an2v0x2_0_b mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1050 diff2_2_xnr2v8x05_0_an diff2_2_in_a mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1051 diff2_2_xnr2v8x05_0_zn diff2_2_in_b diff2_2_xnr2v8x05_0_an mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1052 diff2_2_xnr2v8x05_0_ai diff2_2_xnr2v8x05_0_bn diff2_2_xnr2v8x05_0_zn mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1053 mux_0_gnd diff2_2_xnr2v8x05_0_an diff2_2_xnr2v8x05_0_ai mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1054 diff2_2_xnr2v8x05_0_bn diff2_2_in_b mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1055 diff2_2_an2v0x2_2_a mux_0_a2 mux_0_vdd mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1056 mux_0_vdd mux_0_a2 diff2_2_an2v0x2_2_a mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1057 diff2_2_an2v0x2_2_a mux_0_a2 mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1058 mux_0_gnd mux_0_a2 diff2_2_an2v0x2_2_a mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1059 diff2_2_xor3v1x2_0_cn diff2_2_xor3v1x2_0_zn mux_0_a2 mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1060 mux_0_a2 diff2_2_xor3v1x2_0_zn diff2_2_xor3v1x2_0_cn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1061 diff2_2_xor3v1x2_0_zn diff2_2_xor3v1x2_0_cn mux_0_a2 mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1062 mux_0_a2 diff2_2_xor3v1x2_0_cn diff2_2_xor3v1x2_0_zn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1063 diff2_2_xor3v1x2_0_cn diff2_2_in_c mux_0_vdd mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1064 mux_0_vdd diff2_2_in_c diff2_2_xor3v1x2_0_cn mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1065 diff2_2_xor3v1x2_0_zn diff2_2_xor3v1x2_0_iz mux_0_vdd mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1066 mux_0_vdd diff2_2_xor3v1x2_0_iz diff2_2_xor3v1x2_0_zn mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1067 diff2_2_xor3v1x2_0_iz diff2_2_an2v0x2_1_a diff2_2_xor3v1x2_0_bn mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1068 diff2_2_an2v0x2_1_a diff2_2_xor3v1x2_0_bn diff2_2_xor3v1x2_0_iz mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1069 mux_0_vdd diff2_2_in_a diff2_2_an2v0x2_1_a mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1070 diff2_2_xor3v1x2_0_bn diff2_2_in_b mux_0_vdd mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1071 mux_0_vdd diff2_2_in_b diff2_2_xor3v1x2_0_bn mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1072 diff2_2_xor3v1x2_0_a_11_12# diff2_2_xor3v1x2_0_cn mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1073 mux_0_a2 diff2_2_xor3v1x2_0_zn diff2_2_xor3v1x2_0_a_11_12# mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1074 diff2_2_xor3v1x2_0_a_28_12# diff2_2_xor3v1x2_0_zn mux_0_a2 mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1075 mux_0_gnd diff2_2_xor3v1x2_0_cn diff2_2_xor3v1x2_0_a_28_12# mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1076 diff2_2_xor3v1x2_0_zn diff2_2_xor3v1x2_0_iz mux_0_gnd mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1077 mux_0_a2 diff2_2_in_c diff2_2_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1078 diff2_2_xor3v1x2_0_zn diff2_2_in_c mux_0_a2 mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1079 mux_0_gnd diff2_2_xor3v1x2_0_iz diff2_2_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1080 diff2_2_xor3v1x2_0_cn diff2_2_in_c mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1081 mux_0_gnd diff2_2_in_c diff2_2_xor3v1x2_0_cn mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1082 diff2_2_xor3v1x2_0_a_115_7# diff2_2_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1083 diff2_2_xor3v1x2_0_iz diff2_2_xor3v1x2_0_bn diff2_2_xor3v1x2_0_a_115_7# mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1084 diff2_2_an2v0x2_1_a diff2_2_in_b diff2_2_xor3v1x2_0_iz mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1085 mux_0_gnd diff2_2_in_a diff2_2_an2v0x2_1_a mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1086 diff2_2_xor3v1x2_0_bn diff2_2_in_b mux_0_gnd mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1087 mux_0_vdd diff2_1_an2v0x2_2_zn diff2_2_in_2c mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1088 diff2_1_an2v0x2_2_zn diff2_1_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1089 mux_0_vdd diff2_1_in_2c diff2_1_an2v0x2_2_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1090 mux_0_gnd diff2_1_an2v0x2_2_zn diff2_2_in_2c mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1091 diff2_1_an2v0x2_2_a_24_13# diff2_1_an2v0x2_2_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1092 diff2_1_an2v0x2_2_zn diff2_1_in_2c diff2_1_an2v0x2_2_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1093 diff2_1_xor2v2x2_0_an diff2_1_xor2v2x2_0_bn mux_0_b1 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1094 mux_0_b1 diff2_1_xor2v2x2_0_bn diff2_1_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1095 diff2_1_xor2v2x2_0_bn diff2_1_xor2v2x2_0_an mux_0_b1 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1096 mux_0_b1 diff2_1_xor2v2x2_0_an diff2_1_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1097 diff2_1_xor2v2x2_0_bn diff2_1_in_2c mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1098 mux_0_vdd diff2_1_in_2c diff2_1_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1099 diff2_1_xor2v2x2_0_an diff2_1_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1100 mux_0_vdd diff2_1_an2v0x2_2_a diff2_1_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1101 diff2_1_xor2v2x2_0_a_13_13# diff2_1_xor2v2x2_0_an mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1102 mux_0_b1 diff2_1_xor2v2x2_0_bn diff2_1_xor2v2x2_0_a_13_13# mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1103 diff2_1_xor2v2x2_0_a_30_13# diff2_1_xor2v2x2_0_bn mux_0_b1 mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1104 mux_0_gnd diff2_1_xor2v2x2_0_an diff2_1_xor2v2x2_0_a_30_13# mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1105 diff2_1_xor2v2x2_0_bn diff2_1_in_2c mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1106 mux_0_b1 diff2_1_an2v0x2_2_a diff2_1_xor2v2x2_0_bn mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1107 diff2_1_xor2v2x2_0_an diff2_1_in_2c mux_0_b1 mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1108 mux_0_gnd diff2_1_an2v0x2_2_a diff2_1_xor2v2x2_0_an mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1109 diff2_2_in_c diff2_1_or2v0x3_0_zn mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1110 mux_0_vdd diff2_1_or2v0x3_0_zn diff2_2_in_c mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1111 diff2_1_or2v0x3_0_a_31_39# diff2_1_an2v0x2_1_z mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1112 diff2_1_or2v0x3_0_zn diff2_1_an2v0x2_0_z diff2_1_or2v0x3_0_a_31_39# mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1113 diff2_1_or2v0x3_0_a_48_39# diff2_1_an2v0x2_0_z diff2_1_or2v0x3_0_zn mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1114 mux_0_vdd diff2_1_an2v0x2_1_z diff2_1_or2v0x3_0_a_48_39# mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1115 mux_0_gnd diff2_1_or2v0x3_0_zn diff2_2_in_c mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1116 diff2_1_or2v0x3_0_zn diff2_1_an2v0x2_1_z mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1117 mux_0_gnd diff2_1_an2v0x2_0_z diff2_1_or2v0x3_0_zn mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1118 mux_0_vdd diff2_1_an2v0x2_1_zn diff2_1_an2v0x2_1_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1119 diff2_1_an2v0x2_1_zn diff2_1_an2v0x2_1_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1120 mux_0_vdd diff2_1_in_b diff2_1_an2v0x2_1_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1121 mux_0_gnd diff2_1_an2v0x2_1_zn diff2_1_an2v0x2_1_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1122 diff2_1_an2v0x2_1_a_24_13# diff2_1_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1123 diff2_1_an2v0x2_1_zn diff2_1_in_b diff2_1_an2v0x2_1_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1124 mux_0_vdd diff2_1_an2v0x2_0_zn diff2_1_an2v0x2_0_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1125 diff2_1_an2v0x2_0_zn diff2_1_in_c mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1126 mux_0_vdd diff2_1_an2v0x2_0_b diff2_1_an2v0x2_0_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1127 mux_0_gnd diff2_1_an2v0x2_0_zn diff2_1_an2v0x2_0_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1128 diff2_1_an2v0x2_0_a_24_13# diff2_1_in_c mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1129 diff2_1_an2v0x2_0_zn diff2_1_an2v0x2_0_b diff2_1_an2v0x2_0_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1130 mux_0_vdd diff2_1_xnr2v8x05_0_zn diff2_1_an2v0x2_0_b mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1131 diff2_1_xnr2v8x05_0_an diff2_1_in_a mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1132 diff2_1_xnr2v8x05_0_zn diff2_1_xnr2v8x05_0_bn diff2_1_xnr2v8x05_0_an mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1133 diff2_1_xnr2v8x05_0_ai diff2_1_in_b diff2_1_xnr2v8x05_0_zn mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1134 mux_0_vdd diff2_1_xnr2v8x05_0_an diff2_1_xnr2v8x05_0_ai mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1135 diff2_1_xnr2v8x05_0_bn diff2_1_in_b mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1136 mux_0_gnd diff2_1_xnr2v8x05_0_zn diff2_1_an2v0x2_0_b mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1137 diff2_1_xnr2v8x05_0_an diff2_1_in_a mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1138 diff2_1_xnr2v8x05_0_zn diff2_1_in_b diff2_1_xnr2v8x05_0_an mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1139 diff2_1_xnr2v8x05_0_ai diff2_1_xnr2v8x05_0_bn diff2_1_xnr2v8x05_0_zn mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1140 mux_0_gnd diff2_1_xnr2v8x05_0_an diff2_1_xnr2v8x05_0_ai mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1141 diff2_1_xnr2v8x05_0_bn diff2_1_in_b mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1142 diff2_1_an2v0x2_2_a mux_0_a1 mux_0_vdd mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1143 mux_0_vdd mux_0_a1 diff2_1_an2v0x2_2_a mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1144 diff2_1_an2v0x2_2_a mux_0_a1 mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1145 mux_0_gnd mux_0_a1 diff2_1_an2v0x2_2_a mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1146 diff2_1_xor3v1x2_0_cn diff2_1_xor3v1x2_0_zn mux_0_a1 mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1147 mux_0_a1 diff2_1_xor3v1x2_0_zn diff2_1_xor3v1x2_0_cn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1148 diff2_1_xor3v1x2_0_zn diff2_1_xor3v1x2_0_cn mux_0_a1 mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1149 mux_0_a1 diff2_1_xor3v1x2_0_cn diff2_1_xor3v1x2_0_zn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1150 diff2_1_xor3v1x2_0_cn diff2_1_in_c mux_0_vdd mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1151 mux_0_vdd diff2_1_in_c diff2_1_xor3v1x2_0_cn mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1152 diff2_1_xor3v1x2_0_zn diff2_1_xor3v1x2_0_iz mux_0_vdd mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1153 mux_0_vdd diff2_1_xor3v1x2_0_iz diff2_1_xor3v1x2_0_zn mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1154 diff2_1_xor3v1x2_0_iz diff2_1_an2v0x2_1_a diff2_1_xor3v1x2_0_bn mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1155 diff2_1_an2v0x2_1_a diff2_1_xor3v1x2_0_bn diff2_1_xor3v1x2_0_iz mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1156 mux_0_vdd diff2_1_in_a diff2_1_an2v0x2_1_a mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1157 diff2_1_xor3v1x2_0_bn diff2_1_in_b mux_0_vdd mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1158 mux_0_vdd diff2_1_in_b diff2_1_xor3v1x2_0_bn mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1159 diff2_1_xor3v1x2_0_a_11_12# diff2_1_xor3v1x2_0_cn mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1160 mux_0_a1 diff2_1_xor3v1x2_0_zn diff2_1_xor3v1x2_0_a_11_12# mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1161 diff2_1_xor3v1x2_0_a_28_12# diff2_1_xor3v1x2_0_zn mux_0_a1 mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1162 mux_0_gnd diff2_1_xor3v1x2_0_cn diff2_1_xor3v1x2_0_a_28_12# mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1163 diff2_1_xor3v1x2_0_zn diff2_1_xor3v1x2_0_iz mux_0_gnd mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1164 mux_0_a1 diff2_1_in_c diff2_1_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1165 diff2_1_xor3v1x2_0_zn diff2_1_in_c mux_0_a1 mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1166 mux_0_gnd diff2_1_xor3v1x2_0_iz diff2_1_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1167 diff2_1_xor3v1x2_0_cn diff2_1_in_c mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1168 mux_0_gnd diff2_1_in_c diff2_1_xor3v1x2_0_cn mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1169 diff2_1_xor3v1x2_0_a_115_7# diff2_1_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1170 diff2_1_xor3v1x2_0_iz diff2_1_xor3v1x2_0_bn diff2_1_xor3v1x2_0_a_115_7# mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1171 diff2_1_an2v0x2_1_a diff2_1_in_b diff2_1_xor3v1x2_0_iz mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1172 mux_0_gnd diff2_1_in_a diff2_1_an2v0x2_1_a mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1173 diff2_1_xor3v1x2_0_bn diff2_1_in_b mux_0_gnd mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1174 mux_0_vdd diff2_0_an2v0x2_2_zn diff2_1_in_2c mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1175 diff2_0_an2v0x2_2_zn diff2_0_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1176 mux_0_vdd mux_0_vdd diff2_0_an2v0x2_2_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1177 mux_0_gnd diff2_0_an2v0x2_2_zn diff2_1_in_2c mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1178 diff2_0_an2v0x2_2_a_24_13# diff2_0_an2v0x2_2_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1179 diff2_0_an2v0x2_2_zn mux_0_vdd diff2_0_an2v0x2_2_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1180 diff2_0_xor2v2x2_0_an diff2_0_xor2v2x2_0_bn mux_0_b0 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=398p ps=164u
M1181 mux_0_b0 diff2_0_xor2v2x2_0_bn diff2_0_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1182 diff2_0_xor2v2x2_0_bn diff2_0_xor2v2x2_0_an mux_0_b0 mux_0_vdd pfet w=20u l=2u
+  ad=320p pd=112u as=0p ps=0u
M1183 mux_0_b0 diff2_0_xor2v2x2_0_an diff2_0_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1184 diff2_0_xor2v2x2_0_bn mux_0_vdd mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1185 mux_0_vdd mux_0_vdd diff2_0_xor2v2x2_0_bn mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1186 diff2_0_xor2v2x2_0_an diff2_0_an2v0x2_2_a mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1187 mux_0_vdd diff2_0_an2v0x2_2_a diff2_0_xor2v2x2_0_an mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1188 diff2_0_xor2v2x2_0_a_13_13# diff2_0_xor2v2x2_0_an mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1189 mux_0_b0 diff2_0_xor2v2x2_0_bn diff2_0_xor2v2x2_0_a_13_13# mux_0_gnd nfet w=13u l=2u
+  ad=264p pd=98u as=0p ps=0u
M1190 diff2_0_xor2v2x2_0_a_30_13# diff2_0_xor2v2x2_0_bn mux_0_b0 mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1191 mux_0_gnd diff2_0_xor2v2x2_0_an diff2_0_xor2v2x2_0_a_30_13# mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1192 diff2_0_xor2v2x2_0_bn mux_0_vdd mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1193 mux_0_b0 diff2_0_an2v0x2_2_a diff2_0_xor2v2x2_0_bn mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1194 diff2_0_xor2v2x2_0_an mux_0_vdd mux_0_b0 mux_0_gnd nfet w=20u l=2u
+  ad=130p pd=56u as=0p ps=0u
M1195 mux_0_gnd diff2_0_an2v0x2_2_a diff2_0_xor2v2x2_0_an mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1196 diff2_1_in_c diff2_0_or2v0x3_0_zn mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=160p pd=56u as=0p ps=0u
M1197 mux_0_vdd diff2_0_or2v0x3_0_zn diff2_1_in_c mux_0_vdd pfet w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1198 diff2_0_or2v0x3_0_a_31_39# diff2_0_an2v0x2_1_z mux_0_vdd mux_0_vdd pfet w=20u l=2u
+  ad=100p pd=50u as=0p ps=0u
M1199 diff2_0_or2v0x3_0_zn diff2_0_an2v0x2_0_z diff2_0_or2v0x3_0_a_31_39# mux_0_vdd pfet w=20u l=2u
+  ad=148p pd=56u as=0p ps=0u
M1200 diff2_0_or2v0x3_0_a_48_39# diff2_0_an2v0x2_0_z diff2_0_or2v0x3_0_zn mux_0_vdd pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1201 mux_0_vdd diff2_0_an2v0x2_1_z diff2_0_or2v0x3_0_a_48_39# mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1202 mux_0_gnd diff2_0_or2v0x3_0_zn diff2_1_in_c mux_0_gnd nfet w=20u l=2u
+  ad=0p pd=0u as=126p ps=54u
M1203 diff2_0_or2v0x3_0_zn diff2_0_an2v0x2_1_z mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1204 mux_0_gnd diff2_0_an2v0x2_0_z diff2_0_or2v0x3_0_zn mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1205 mux_0_vdd diff2_0_an2v0x2_1_zn diff2_0_an2v0x2_1_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1206 diff2_0_an2v0x2_1_zn diff2_0_an2v0x2_1_a mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1207 mux_0_vdd diff2_0_in_b diff2_0_an2v0x2_1_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1208 mux_0_gnd diff2_0_an2v0x2_1_zn diff2_0_an2v0x2_1_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1209 diff2_0_an2v0x2_1_a_24_13# diff2_0_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1210 diff2_0_an2v0x2_1_zn diff2_0_in_b diff2_0_an2v0x2_1_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1211 mux_0_vdd diff2_0_an2v0x2_0_zn diff2_0_an2v0x2_0_z mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=166p ps=70u
M1212 diff2_0_an2v0x2_0_zn mux_0_gnd mux_0_vdd mux_0_vdd pfet w=19u l=2u
+  ad=152p pd=54u as=0p ps=0u
M1213 mux_0_vdd diff2_0_an2v0x2_0_b diff2_0_an2v0x2_0_zn mux_0_vdd pfet w=19u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1214 mux_0_gnd diff2_0_an2v0x2_0_zn diff2_0_an2v0x2_0_z mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=98p ps=42u
M1215 diff2_0_an2v0x2_0_a_24_13# mux_0_gnd mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1216 diff2_0_an2v0x2_0_zn diff2_0_an2v0x2_0_b diff2_0_an2v0x2_0_a_24_13# mux_0_gnd nfet w=13u l=2u
+  ad=77p pd=40u as=0p ps=0u
M1217 mux_0_vdd diff2_0_xnr2v8x05_0_zn diff2_0_an2v0x2_0_b mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=72p ps=38u
M1218 diff2_0_xnr2v8x05_0_an diff2_0_in_a mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1219 diff2_0_xnr2v8x05_0_zn diff2_0_xnr2v8x05_0_bn diff2_0_xnr2v8x05_0_an mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1220 diff2_0_xnr2v8x05_0_ai diff2_0_in_b diff2_0_xnr2v8x05_0_zn mux_0_vdd pfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1221 mux_0_vdd diff2_0_xnr2v8x05_0_an diff2_0_xnr2v8x05_0_ai mux_0_vdd pfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1222 diff2_0_xnr2v8x05_0_bn diff2_0_in_b mux_0_vdd mux_0_vdd pfet w=12u l=2u
+  ad=72p pd=38u as=0p ps=0u
M1223 mux_0_gnd diff2_0_xnr2v8x05_0_zn diff2_0_an2v0x2_0_b mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=42p ps=26u
M1224 diff2_0_xnr2v8x05_0_an diff2_0_in_a mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1225 diff2_0_xnr2v8x05_0_zn diff2_0_in_b diff2_0_xnr2v8x05_0_an mux_0_gnd nfet w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1226 diff2_0_xnr2v8x05_0_ai diff2_0_xnr2v8x05_0_bn diff2_0_xnr2v8x05_0_zn mux_0_gnd nfet w=6u l=2u
+  ad=57p pd=32u as=0p ps=0u
M1227 mux_0_gnd diff2_0_xnr2v8x05_0_an diff2_0_xnr2v8x05_0_ai mux_0_gnd nfet w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1228 diff2_0_xnr2v8x05_0_bn diff2_0_in_b mux_0_gnd mux_0_gnd nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1229 diff2_0_an2v0x2_2_a mux_0_a0 mux_0_vdd mux_0_vdd pfet w=24u l=2u
+  ad=168p pd=64u as=0p ps=0u
M1230 mux_0_vdd mux_0_a0 diff2_0_an2v0x2_2_a mux_0_vdd pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1231 diff2_0_an2v0x2_2_a mux_0_a0 mux_0_gnd mux_0_gnd nfet w=10u l=2u
+  ad=80p pd=36u as=0p ps=0u
M1232 mux_0_gnd mux_0_a0 diff2_0_an2v0x2_2_a mux_0_gnd nfet w=10u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1233 diff2_0_xor3v1x2_0_cn diff2_0_xor3v1x2_0_zn mux_0_a0 mux_0_vdd pfet w=27u l=2u
+  ad=424p pd=138u as=530p ps=208u
M1234 mux_0_a0 diff2_0_xor3v1x2_0_zn diff2_0_xor3v1x2_0_cn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1235 diff2_0_xor3v1x2_0_zn diff2_0_xor3v1x2_0_cn mux_0_a0 mux_0_vdd pfet w=27u l=2u
+  ad=440p pd=142u as=0p ps=0u
M1236 mux_0_a0 diff2_0_xor3v1x2_0_cn diff2_0_xor3v1x2_0_zn mux_0_vdd pfet w=27u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1237 diff2_0_xor3v1x2_0_cn mux_0_gnd mux_0_vdd mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1238 mux_0_vdd mux_0_gnd diff2_0_xor3v1x2_0_cn mux_0_vdd pfet w=26u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1239 diff2_0_xor3v1x2_0_zn diff2_0_xor3v1x2_0_iz mux_0_vdd mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1240 mux_0_vdd diff2_0_xor3v1x2_0_iz diff2_0_xor3v1x2_0_zn mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1241 diff2_0_xor3v1x2_0_iz diff2_0_an2v0x2_1_a diff2_0_xor3v1x2_0_bn mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=272p ps=122u
M1242 diff2_0_an2v0x2_1_a diff2_0_xor3v1x2_0_bn diff2_0_xor3v1x2_0_iz mux_0_vdd pfet w=28u l=2u
+  ad=224p pd=72u as=0p ps=0u
M1243 mux_0_vdd diff2_0_in_a diff2_0_an2v0x2_1_a mux_0_vdd pfet w=28u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1244 diff2_0_xor3v1x2_0_bn diff2_0_in_b mux_0_vdd mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1245 mux_0_vdd diff2_0_in_b diff2_0_xor3v1x2_0_bn mux_0_vdd pfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1246 diff2_0_xor3v1x2_0_a_11_12# diff2_0_xor3v1x2_0_cn mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1247 mux_0_a0 diff2_0_xor3v1x2_0_zn diff2_0_xor3v1x2_0_a_11_12# mux_0_gnd nfet w=12u l=2u
+  ad=208p pd=84u as=0p ps=0u
M1248 diff2_0_xor3v1x2_0_a_28_12# diff2_0_xor3v1x2_0_zn mux_0_a0 mux_0_gnd nfet w=12u l=2u
+  ad=60p pd=34u as=0p ps=0u
M1249 mux_0_gnd diff2_0_xor3v1x2_0_cn diff2_0_xor3v1x2_0_a_28_12# mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1250 diff2_0_xor3v1x2_0_zn diff2_0_xor3v1x2_0_iz mux_0_gnd mux_0_gnd nfet w=14u l=2u
+  ad=224p pd=88u as=0p ps=0u
M1251 mux_0_a0 mux_0_gnd diff2_0_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1252 diff2_0_xor3v1x2_0_zn mux_0_gnd mux_0_a0 mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1253 mux_0_gnd diff2_0_xor3v1x2_0_iz diff2_0_xor3v1x2_0_zn mux_0_gnd nfet w=14u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1254 diff2_0_xor3v1x2_0_cn mux_0_gnd mux_0_gnd mux_0_gnd nfet w=12u l=2u
+  ad=96p pd=40u as=0p ps=0u
M1255 mux_0_gnd mux_0_gnd diff2_0_xor3v1x2_0_cn mux_0_gnd nfet w=12u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1256 diff2_0_xor3v1x2_0_a_115_7# diff2_0_an2v0x2_1_a mux_0_gnd mux_0_gnd nfet w=13u l=2u
+  ad=65p pd=36u as=0p ps=0u
M1257 diff2_0_xor3v1x2_0_iz diff2_0_xor3v1x2_0_bn diff2_0_xor3v1x2_0_a_115_7# mux_0_gnd nfet w=13u l=2u
+  ad=104p pd=42u as=0p ps=0u
M1258 diff2_0_an2v0x2_1_a diff2_0_in_b diff2_0_xor3v1x2_0_iz mux_0_gnd nfet w=13u l=2u
+  ad=114p pd=52u as=0p ps=0u
M1259 mux_0_gnd diff2_0_in_a diff2_0_an2v0x2_1_a mux_0_gnd nfet w=13u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1260 diff2_0_xor3v1x2_0_bn diff2_0_in_b mux_0_gnd mux_0_gnd nfet w=11u l=2u
+  ad=67p pd=36u as=0p ps=0u
M1261 mux_0_vdd mux_0_mxn2v0x1_2_zn mux_0_o2 mux_0_mxn2v0x1_1_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1262 mux_0_mxn2v0x1_2_a_21_50# mux_0_a2 mux_0_vdd mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1263 mux_0_mxn2v0x1_2_zn mux_0_s mux_0_mxn2v0x1_2_a_21_50# mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1264 mux_0_mxn2v0x1_2_a_38_50# mux_0_mxn2v0x1_2_sn mux_0_mxn2v0x1_2_zn mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1265 mux_0_vdd mux_0_b2 mux_0_mxn2v0x1_2_a_38_50# mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1266 mux_0_mxn2v0x1_2_sn mux_0_s mux_0_vdd mux_0_mxn2v0x1_1_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1267 mux_0_gnd mux_0_mxn2v0x1_2_zn mux_0_o2 mux_0_mxn2v0x1_2_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1268 mux_0_mxn2v0x1_2_a_21_12# mux_0_a2 mux_0_gnd mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1269 mux_0_mxn2v0x1_2_zn mux_0_mxn2v0x1_2_sn mux_0_mxn2v0x1_2_a_21_12# mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1270 mux_0_mxn2v0x1_2_a_38_12# mux_0_s mux_0_mxn2v0x1_2_zn mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1271 mux_0_gnd mux_0_b2 mux_0_mxn2v0x1_2_a_38_12# mux_0_mxn2v0x1_2_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1272 mux_0_mxn2v0x1_2_sn mux_0_s mux_0_gnd mux_0_mxn2v0x1_2_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1273 mux_0_vdd mux_0_mxn2v0x1_1_zn mux_0_o1 mux_0_mxn2v0x1_1_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1274 mux_0_mxn2v0x1_1_a_21_50# mux_0_a1 mux_0_vdd mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1275 mux_0_mxn2v0x1_1_zn mux_0_s mux_0_mxn2v0x1_1_a_21_50# mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1276 mux_0_mxn2v0x1_1_a_38_50# mux_0_mxn2v0x1_1_sn mux_0_mxn2v0x1_1_zn mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1277 mux_0_vdd mux_0_b1 mux_0_mxn2v0x1_1_a_38_50# mux_0_mxn2v0x1_1_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1278 mux_0_mxn2v0x1_1_sn mux_0_s mux_0_vdd mux_0_mxn2v0x1_1_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1279 mux_0_gnd mux_0_mxn2v0x1_1_zn mux_0_o1 mux_0_mxn2v0x1_0_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1280 mux_0_mxn2v0x1_1_a_21_12# mux_0_a1 mux_0_gnd mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1281 mux_0_mxn2v0x1_1_zn mux_0_mxn2v0x1_1_sn mux_0_mxn2v0x1_1_a_21_12# mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1282 mux_0_mxn2v0x1_1_a_38_12# mux_0_s mux_0_mxn2v0x1_1_zn mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1283 mux_0_gnd mux_0_b1 mux_0_mxn2v0x1_1_a_38_12# mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1284 mux_0_mxn2v0x1_1_sn mux_0_s mux_0_gnd mux_0_mxn2v0x1_0_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1285 mux_0_vdd mux_0_mxn2v0x1_0_zn mux_0_o0 mux_0_mxn2v0x1_0_w_n4_32# pfet w=18u l=2u
+  ad=0p pd=0u as=102p ps=50u
M1286 mux_0_mxn2v0x1_0_a_21_50# mux_0_a0 mux_0_vdd mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1287 mux_0_mxn2v0x1_0_zn mux_0_s mux_0_mxn2v0x1_0_a_21_50# mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=128p pd=48u as=0p ps=0u
M1288 mux_0_mxn2v0x1_0_a_38_50# mux_0_mxn2v0x1_0_sn mux_0_mxn2v0x1_0_zn mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=80p pd=42u as=0p ps=0u
M1289 mux_0_vdd mux_0_b0 mux_0_mxn2v0x1_0_a_38_50# mux_0_mxn2v0x1_0_w_n4_32# pfet w=16u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1290 mux_0_mxn2v0x1_0_sn mux_0_s mux_0_vdd mux_0_mxn2v0x1_0_w_n4_32# pfet w=8u l=2u
+  ad=52p pd=30u as=0p ps=0u
M1291 mux_0_gnd mux_0_mxn2v0x1_0_zn mux_0_o0 mux_0_mxn2v0x1_0_w_n4_n4# nfet w=9u l=2u
+  ad=0p pd=0u as=57p ps=32u
M1292 mux_0_mxn2v0x1_0_a_21_12# mux_0_a0 mux_0_gnd mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1293 mux_0_mxn2v0x1_0_zn mux_0_mxn2v0x1_0_sn mux_0_mxn2v0x1_0_a_21_12# mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=64p pd=32u as=0p ps=0u
M1294 mux_0_mxn2v0x1_0_a_38_12# mux_0_s mux_0_mxn2v0x1_0_zn mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1295 mux_0_gnd mux_0_b0 mux_0_mxn2v0x1_0_a_38_12# mux_0_mxn2v0x1_0_w_n4_n4# nfet w=8u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1296 mux_0_mxn2v0x1_0_sn mux_0_s mux_0_gnd mux_0_mxn2v0x1_0_w_n4_n4# nfet w=6u l=2u
+  ad=42p pd=26u as=0p ps=0u
C0 mux_0_vdd diff2_0_an2v0x2_0_z 24.6fF
C1 diff2_0_xor3v1x2_0_bn mux_0_gnd 9.1fF
C2 diff2_1_xor3v1x2_0_zn diff2_1_in_b 4.3fF
C3 diff2_2_xor3v1x2_0_iz mux_0_gnd 24.9fF
C4 diff2_0_an2v0x2_1_a diff2_0_in_b 2.0fF
C5 mux_0_vdd diff2_1_xor3v1x2_0_cn 31.6fF
C6 diff2_0_xor3v1x2_0_zn mux_0_gnd 13.9fF
C7 diff2_2_xnr2v8x05_0_bn mux_0_vdd 14.4fF
C8 diff2_2_an2v0x2_1_zn mux_0_gnd 8.9fF
C9 diff2_2_an2v0x2_0_zn mux_0_vdd 8.8fF
C10 diff2_1_an2v0x2_0_z mux_0_gnd 12.8fF
C11 mux_0_vdd diff2_0_xor2v2x2_0_an 27.4fF
C12 diff2_2_an2v0x2_1_a mux_0_vdd 12.4fF
C13 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_a1 4.8fF
C14 mux_0_mxn2v0x1_1_w_n4_32# mux_0_o2 6.3fF
C15 diff2_0_an2v0x2_0_z mux_0_gnd 12.8fF
C16 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_gnd 76.0fF
C17 diff2_1_xor3v1x2_0_cn mux_0_a1 4.1fF
C18 diff2_1_an2v0x2_1_z mux_0_vdd 17.7fF
C19 diff2_1_xor2v2x2_0_an mux_0_b1 3.9fF
C20 diff2_1_xor3v1x2_0_cn mux_0_gnd 18.8fF
C21 diff2_0_xor3v1x2_0_iz diff2_0_xor3v1x2_0_bn 2.4fF
C22 mux_0_vdd diff2_0_xor2v2x2_0_bn 18.7fF
C23 diff2_2_xnr2v8x05_0_zn diff2_2_in_c 3.1fF
C24 diff2_2_xnr2v8x05_0_bn mux_0_gnd 6.7fF
C25 mux_0_vdd diff2_0_an2v0x2_1_zn 8.8fF
C26 mux_0_mxn2v0x1_0_w_n4_32# mux_0_mxn2v0x1_0_sn 9.3fF
C27 mux_0_vdd diff2_0_in_a 24.6fF
C28 diff2_2_an2v0x2_0_zn diff2_2_in_a 2.2fF
C29 mux_0_a0 mux_0_mxn2v0x1_0_w_n4_32# 11.6fF
C30 mux_0_vdd diff2_1_an2v0x2_1_a 12.4fF
C31 diff2_0_an2v0x2_2_a diff2_0_xor3v1x2_0_cn 2.3fF
C32 mux_0_vdd diff2_0_xor3v1x2_0_cn 31.6fF
C33 diff2_2_an2v0x2_0_zn mux_0_gnd 8.9fF
C34 diff2_0_xor2v2x2_0_an mux_0_gnd 21.6fF
C35 mux_0_vdd diff2_1_xnr2v8x05_0_bn 14.4fF
C36 diff2_2_an2v0x2_1_a mux_0_gnd 19.1fF
C37 mux_0_vdd diff2_0_an2v0x2_1_a 12.4fF
C38 mux_0_vdd diff2_1_an2v0x2_0_zn 8.8fF
C39 diff2_1_an2v0x2_1_z mux_0_gnd 10.2fF
C40 diff2_2_or2v0x3_0_zn mux_0_vdd 12.7fF
C41 diff2_0_xor2v2x2_0_bn mux_0_gnd 11.2fF
C42 mux_0_vdd diff2_0_an2v0x2_2_zn 10.3fF
C43 mux_0_vdd diff2_0_an2v0x2_0_zn 8.8fF
C44 diff2_0_an2v0x2_1_zn mux_0_gnd 8.9fF
C45 mux_0_a0 diff2_0_xor3v1x2_0_zn 4.6fF
C46 diff2_1_or2v0x3_0_zn mux_0_vdd 12.7fF
C47 diff2_0_in_a mux_0_gnd 26.8fF
C48 diff2_1_an2v0x2_1_a mux_0_gnd 19.1fF
C49 mux_0_vdd diff2_1_in_c 39.6fF
C50 diff2_0_xor3v1x2_0_cn mux_0_gnd 19.1fF
C51 mux_0_vdd diff2_0_in_b 50.3fF
C52 mux_0_vdd diff2_2_xor3v1x2_0_bn 15.4fF
C53 diff2_1_xnr2v8x05_0_bn mux_0_gnd 6.7fF
C54 diff2_2_an2v0x2_1_a diff2_2_in_b 2.0fF
C55 mux_0_mxn2v0x1_1_w_n4_32# mux_0_b2 6.6fF
C56 mux_0_vdd mux_0_mxn2v0x1_1_w_n4_32# 59.4fF
C57 diff2_0_an2v0x2_1_a mux_0_gnd 19.1fF
C58 mux_0_vdd mux_0_b0 26.2fF
C59 mux_0_mxn2v0x1_0_w_n4_32# mux_0_o0 5.2fF
C60 mux_0_vdd diff2_2_xor3v1x2_0_zn 18.9fF
C61 mux_0_vdd diff2_1_xnr2v8x05_0_an 9.9fF
C62 mux_0_vdd diff2_1_xor3v1x2_0_bn 15.4fF
C63 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_mxn2v0x1_0_sn 9.2fF
C64 diff2_1_an2v0x2_0_zn mux_0_gnd 8.9fF
C65 mux_0_a0 mux_0_mxn2v0x1_0_w_n4_n4# 4.8fF
C66 mux_0_mxn2v0x1_0_w_n4_32# mux_0_mxn2v0x1_0_zn 9.3fF
C67 diff2_2_or2v0x3_0_zn mux_0_gnd 9.0fF
C68 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_mxn2v0x1_1_sn 9.2fF
C69 mux_0_vdd diff2_0_xnr2v8x05_0_bn 14.4fF
C70 diff2_1_an2v0x2_0_zn diff2_1_in_a 2.2fF
C71 diff2_0_an2v0x2_2_zn mux_0_gnd 8.9fF
C72 diff2_2_an2v0x2_1_z mux_0_vdd 17.7fF
C73 diff2_0_an2v0x2_0_zn mux_0_gnd 10.8fF
C74 diff2_0_an2v0x2_1_z mux_0_vdd 17.7fF
C75 diff2_1_or2v0x3_0_zn mux_0_gnd 9.0fF
C76 mux_0_mxn2v0x1_1_w_n4_32# mux_0_a1 13.4fF
C77 diff2_1_in_c mux_0_gnd 33.4fF
C78 diff2_2_an2v0x2_2_zn mux_0_vdd 8.8fF
C79 diff2_0_in_b mux_0_gnd 56.4fF
C80 diff2_2_xor3v1x2_0_bn mux_0_gnd 9.1fF
C81 mux_0_mxn2v0x1_0_w_n4_32# mux_0_s 18.7fF
C82 diff2_1_an2v0x2_1_a diff2_1_in_b 2.0fF
C83 mux_0_b0 mux_0_gnd 10.9fF
C84 diff2_2_xor3v1x2_0_zn diff2_2_xor3v1x2_0_cn 4.5fF
C85 diff2_2_xor3v1x2_0_zn mux_0_gnd 11.9fF
C86 diff2_1_xnr2v8x05_0_an mux_0_gnd 5.5fF
C87 mux_0_vdd diff2_1_an2v0x2_2_a 59.6fF
C88 diff2_1_xor3v1x2_0_bn mux_0_gnd 9.1fF
C89 mux_0_o1 mux_0_mxn2v0x1_0_w_n4_n4# 2.3fF
C90 mux_0_mxn2v0x1_2_w_n4_n4# mux_0_o2 2.3fF
C91 diff2_0_xnr2v8x05_0_bn mux_0_gnd 7.5fF
C92 mux_0_vdd diff2_0_an2v0x2_2_a 61.1fF
C93 mux_0_vdd mux_0_b2 13.6fF
C94 diff2_2_an2v0x2_1_z mux_0_gnd 10.2fF
C95 mux_0_vdd diff2_0_xnr2v8x05_0_an 9.9fF
C96 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_o0 2.3fF
C97 diff2_0_an2v0x2_1_z mux_0_gnd 10.2fF
C98 diff2_2_an2v0x2_0_z mux_0_vdd 24.6fF
C99 diff2_2_an2v0x2_2_zn mux_0_gnd 8.9fF
C100 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_mxn2v0x1_0_zn 8.9fF
C101 diff2_2_xor3v1x2_0_bn diff2_2_in_b 2.6fF
C102 mux_0_a0 diff2_0_xor3v1x2_0_cn 4.1fF
C103 mux_0_mxn2v0x1_1_w_n4_32# mux_0_mxn2v0x1_2_zn 9.3fF
C104 diff2_2_xor3v1x2_0_zn diff2_2_in_b 4.3fF
C105 diff2_1_an2v0x2_2_a mux_0_gnd 25.3fF
C106 diff2_1_xnr2v8x05_0_zn diff2_1_in_c 3.1fF
C107 mux_0_vdd mux_0_a1 38.3fF
C108 mux_0_vdd diff2_2_in_a 24.6fF
C109 diff2_0_an2v0x2_2_a mux_0_gnd 25.3fF
C110 mux_0_vdd diff2_2_xor3v1x2_0_cn 31.6fF
C111 mux_0_vdd mux_0_gnd 45.8fF
C112 diff2_1_xor3v1x2_0_bn diff2_1_in_b 2.6fF
C113 mux_0_b2 mux_0_gnd 15.7fF
C114 mux_0_vdd diff2_1_in_a 24.6fF
C115 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_s 30.3fF
C116 diff2_0_xnr2v8x05_0_an mux_0_gnd 6.8fF
C117 mux_0_vdd diff2_1_xor2v2x2_0_bn 17.7fF
C118 diff2_2_an2v0x2_0_z mux_0_gnd 12.8fF
C119 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_b1 10.2fF
C120 diff2_1_xor3v1x2_0_zn diff2_1_xor3v1x2_0_cn 4.5fF
C121 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_mxn2v0x1_1_zn 8.9fF
C122 diff2_2_xor2v2x2_0_bn mux_0_vdd 17.7fF
C123 diff2_2_xor2v2x2_0_bn mux_0_b2 2.7fF
C124 mux_0_vdd diff2_0_an2v0x2_0_b 20.5fF
C125 mux_0_vdd diff2_0_or2v0x3_0_zn 12.7fF
C126 mux_0_mxn2v0x1_1_w_n4_32# mux_0_mxn2v0x1_1_sn 9.3fF
C127 mux_0_mxn2v0x1_2_w_n4_n4# mux_0_b2 8.7fF
C128 diff2_2_in_2c mux_0_vdd 33.2fF
C129 diff2_2_in_a mux_0_gnd 26.6fF
C130 mux_0_gnd mux_0_a1 14.9fF
C131 diff2_2_xnr2v8x05_0_an mux_0_vdd 9.9fF
C132 diff2_2_xor3v1x2_0_cn mux_0_gnd 18.8fF
C133 mux_0_vdd diff2_2_in_b 50.3fF
C134 mux_0_mxn2v0x1_2_zn mux_0_b2 2.7fF
C135 diff2_1_in_a mux_0_gnd 26.6fF
C136 mux_0_vdd diff2_0_xor3v1x2_0_iz 15.8fF
C137 mux_0_vdd diff2_1_an2v0x2_1_zn 8.8fF
C138 diff2_1_xor2v2x2_0_bn mux_0_gnd 11.2fF
C139 mux_0_vdd diff2_1_in_b 50.3fF
C140 mux_0_vdd diff2_1_xnr2v8x05_0_zn 4.4fF
C141 mux_0_vdd diff2_1_an2v0x2_0_b 20.5fF
C142 diff2_2_xor2v2x2_0_bn mux_0_gnd 11.2fF
C143 diff2_0_an2v0x2_0_b mux_0_gnd 7.3fF
C144 mux_0_o1 mux_0_mxn2v0x1_1_w_n4_32# 5.0fF
C145 diff2_0_or2v0x3_0_zn mux_0_gnd 9.0fF
C146 mux_0_mxn2v0x1_2_w_n4_n4# mux_0_gnd 25.5fF
C147 diff2_2_xor2v2x2_0_an mux_0_b2 3.9fF
C148 diff2_2_xor2v2x2_0_an mux_0_vdd 25.5fF
C149 diff2_2_in_2c mux_0_gnd 16.8fF
C150 diff2_2_an2v0x2_2_z mux_0_vdd 2.4fF
C151 diff2_2_xnr2v8x05_0_an mux_0_gnd 5.5fF
C152 diff2_2_in_b mux_0_gnd 56.1fF
C153 diff2_0_xor3v1x2_0_iz mux_0_gnd 25.5fF
C154 mux_0_a0 mux_0_vdd 35.5fF
C155 diff2_1_an2v0x2_1_zn mux_0_gnd 8.9fF
C156 mux_0_a2 mux_0_mxn2v0x1_1_w_n4_32# 11.6fF
C157 diff2_1_in_b mux_0_gnd 56.1fF
C158 mux_0_b0 mux_0_mxn2v0x1_0_zn 2.7fF
C159 diff2_1_xor2v2x2_0_an mux_0_vdd 25.5fF
C160 mux_0_a2 diff2_2_xor3v1x2_0_zn 4.6fF
C161 diff2_1_xnr2v8x05_0_zn mux_0_gnd 11.9fF
C162 diff2_2_an2v0x2_0_b mux_0_vdd 20.5fF
C163 diff2_1_an2v0x2_0_b mux_0_gnd 5.9fF
C164 diff2_2_xor2v2x2_0_an mux_0_gnd 21.6fF
C165 mux_0_vdd diff2_0_xnr2v8x05_0_zn 4.4fF
C166 mux_0_mxn2v0x1_2_zn mux_0_mxn2v0x1_2_w_n4_n4# 8.9fF
C167 mux_0_mxn2v0x1_1_w_n4_32# mux_0_mxn2v0x1_2_sn 9.3fF
C168 mux_0_mxn2v0x1_1_w_n4_32# mux_0_s 36.4fF
C169 diff2_2_an2v0x2_2_z mux_0_gnd 2.5fF
C170 mux_0_mxn2v0x1_1_w_n4_32# mux_0_b1 6.6fF
C171 mux_0_a0 mux_0_gnd 14.9fF
C172 diff2_1_xor2v2x2_0_an mux_0_gnd 21.6fF
C173 diff2_2_xor2v2x2_0_bn diff2_2_xor2v2x2_0_an 3.3fF
C174 mux_0_mxn2v0x1_1_w_n4_32# mux_0_mxn2v0x1_1_zn 9.3fF
C175 diff2_0_xor3v1x2_0_zn diff2_0_xor3v1x2_0_cn 4.5fF
C176 diff2_1_xor2v2x2_0_an diff2_1_xor2v2x2_0_bn 3.3fF
C177 diff2_2_xnr2v8x05_0_zn mux_0_vdd 4.4fF
C178 diff2_2_an2v0x2_0_b mux_0_gnd 5.9fF
C179 mux_0_vdd diff2_2_in_c 40.7fF
C180 mux_0_a2 mux_0_vdd 36.6fF
C181 mux_0_mxn2v0x1_0_w_n4_32# mux_0_b0 6.6fF
C182 diff2_1_xor3v1x2_0_iz diff2_1_xor3v1x2_0_bn 2.4fF
C183 mux_0_vdd diff2_2_an2v0x2_2_a 59.6fF
C184 diff2_0_xnr2v8x05_0_zn mux_0_gnd 15.0fF
C185 diff2_1_an2v0x2_2_zn mux_0_vdd 8.8fF
C186 diff2_0_xor3v1x2_0_bn diff2_0_in_b 2.6fF
C187 diff2_2_xor3v1x2_0_iz diff2_2_xor3v1x2_0_bn 2.4fF
C188 mux_0_vdd mux_0_s 7.9fF
C189 diff2_0_xor3v1x2_0_zn diff2_0_in_b 4.3fF
C190 diff2_0_xor2v2x2_0_bn diff2_0_xor2v2x2_0_an 3.3fF
C191 diff2_2_xnr2v8x05_0_zn mux_0_gnd 11.9fF
C192 mux_0_vdd mux_0_b1 13.2fF
C193 diff2_2_in_c mux_0_gnd 33.4fF
C194 mux_0_vdd diff2_1_xor3v1x2_0_zn 18.9fF
C195 mux_0_a2 diff2_2_xor3v1x2_0_cn 4.1fF
C196 mux_0_a2 mux_0_gnd 14.9fF
C197 diff2_2_an2v0x2_2_a diff2_2_xor3v1x2_0_cn 2.3fF
C198 diff2_2_an2v0x2_2_a mux_0_gnd 25.3fF
C199 diff2_1_in_2c mux_0_vdd 34.0fF
C200 diff2_1_an2v0x2_2_zn mux_0_gnd 8.9fF
C201 mux_0_vdd diff2_1_xor3v1x2_0_iz 15.8fF
C202 mux_0_vdd mux_0_mxn2v0x1_0_w_n4_32# 21.1fF
C203 mux_0_mxn2v0x1_0_w_n4_n4# mux_0_b0 8.7fF
C204 mux_0_gnd mux_0_s 8.3fF
C205 mux_0_a2 mux_0_mxn2v0x1_2_w_n4_n4# 4.8fF
C206 diff2_1_xor3v1x2_0_zn mux_0_a1 4.6fF
C207 mux_0_gnd mux_0_b1 19.6fF
C208 diff2_1_xor3v1x2_0_zn mux_0_gnd 11.9fF
C209 diff2_1_xor2v2x2_0_bn mux_0_b1 2.7fF
C210 mux_0_vdd diff2_0_xor3v1x2_0_bn 15.4fF
C211 diff2_1_in_2c mux_0_gnd 17.5fF
C212 mux_0_vdd diff2_2_xor3v1x2_0_iz 15.8fF
C213 diff2_1_xor3v1x2_0_iz mux_0_gnd 24.9fF
C214 mux_0_vdd diff2_0_xor3v1x2_0_zn 18.9fF
C215 diff2_0_xor2v2x2_0_an mux_0_b0 3.9fF
C216 mux_0_mxn2v0x1_2_w_n4_n4# mux_0_mxn2v0x1_2_sn 9.2fF
C217 mux_0_mxn2v0x1_2_w_n4_n4# mux_0_s 15.2fF
C218 diff2_2_an2v0x2_1_zn mux_0_vdd 8.8fF
C219 diff2_0_an2v0x2_0_zn diff2_0_in_a 2.2fF
C220 mux_0_vdd diff2_1_an2v0x2_0_z 24.6fF
C221 mux_0_o0 mux_0_mxn2v0x1_0_sn 4.3fF
C222 diff2_0_xor2v2x2_0_bn mux_0_b0 2.7fF
C223 mux_0_a0 mux_0_o0 2.3fF
C224 diff2_1_an2v0x2_2_a diff2_1_xor3v1x2_0_cn 2.3fF
C225 mux_0_b0 0 29.8fF
C226 mux_0_s 0 40.5fF
C227 mux_0_a0 0 54.7fF
C228 mux_0_gnd 0 220.8fF
C229 mux_0_o1 0 2.4fF
C230 mux_0_b1 0 25.4fF
C231 mux_0_a1 0 21.5fF
C232 mux_0_b2 0 30.1fF
C233 mux_0_a2 0 20.1fF
C234 diff2_0_in_a 0 4.4fF
C235 diff2_0_an2v0x2_0_b 0 2.9fF
C236 diff2_1_in_c 0 37.1fF
C237 diff2_0_an2v0x2_0_z 0 5.0fF
C238 diff2_1_in_a 0 4.4fF
C239 diff2_1_an2v0x2_0_b 0 2.9fF
C240 diff2_2_in_c 0 37.4fF
C241 diff2_1_an2v0x2_0_z 0 5.0fF
C242 diff2_1_in_2c 0 29.6fF
C243 diff2_2_in_a 0 4.4fF
C244 mux_0_vdd 0 146.5fF
C245 diff2_2_an2v0x2_0_b 0 2.9fF
C246 diff2_2_an2v0x2_0_z 0 5.0fF
C247 diff2_2_in_2c 0 35.3fF

v_ss mux_0_gnd 0 0
v_dd mux_0_vdd 0 5

v_a1 diff2_0_in_a 0 DC 1 PULSE(0 5 0 0 0 20ns 40ns )
v_a2 diff2_1_in_a 0 DC 1 PULSE(0 5 0 0 0 20ns 40ns )
v_a3 diff2_2_in_a 0 DC 1 PULSE(0 5 0 0 0 20ns 40ns )
v_b1 diff2_0_in_b 0 DC 1 PULSE(0 5 0 0 0 40ns 80ns )
v_b2 diff2_1_in_b 0 DC 1 PULSE(0 5 0 0 0 40ns 80ns )
v_b3 diff2_2_in_b 0 DC 1 PULSE(0 5 0 0 0 40ns 80ns )

.tran 0.01ns 200ns 

.control
run 
setplot tran1
plot (mux_0_o0) (mux_0_o1 + 5) (mux_0_o2 + 10)
.endc 

.end