* Sat Apr  9 18:55:28 CEST 2005
.subckt xaon21v0x3 a1 a2 b vdd vss z 
*SPICE circuit <xaon21v0x3> from XCircuit v3.20

m1 an a1 vdd vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m2 n2 a1 vss vss n w=58u l=2u ad='58u*5u+12p' as='58u*5u+12p' pd='58u*2+14u' ps='58u*2+14u'
m3 an a2 n2 vss n w=58u l=2u ad='58u*5u+12p' as='58u*5u+12p' pd='58u*2+14u' ps='58u*2+14u'
m4 bn b vss vss n w=37u l=2u ad='37u*5u+12p' as='37u*5u+12p' pd='37u*2+14u' ps='37u*2+14u'
m5 z bn n1 vss n w=37u l=2u ad='37u*5u+12p' as='37u*5u+12p' pd='37u*2+14u' ps='37u*2+14u'
m6 z b an vss n w=40u l=2u ad='40u*5u+12p' as='40u*5u+12p' pd='40u*2+14u' ps='40u*2+14u'
m7 z bn an vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m8 n1 an vss vss n w=37u l=2u ad='37u*5u+12p' as='37u*5u+12p' pd='37u*2+14u' ps='37u*2+14u'
m9 an a2 vdd vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m10 bn b vdd vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m11 z an bn vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
.ends
