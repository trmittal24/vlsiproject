* Tue Apr  3 09:40:29 CEST 2007
.subckt oai21v0x8 a1 a2 b vdd vss z
*SPICE circuit <oai21v0x8> from XCircuit v3.4 rev 26

m1 n2 a1 vdd vdd p w=217u l=2.3636u ad='217u*5u+12p' as='217u*5u+12p' pd='217u*2+14u' ps='217u*2+14u'
m2 z b vdd vdd p w=112u l=2.3636u ad='112u*5u+12p' as='112u*5u+12p' pd='112u*2+14u' ps='112u*2+14u'
m3 n1 a2 vss vss n w=96u l=2.3636u ad='96u*5u+12p' as='96u*5u+12p' pd='96u*2+14u' ps='96u*2+14u'
m4 n1 a1 vss vss n w=96u l=2.3636u ad='96u*5u+12p' as='96u*5u+12p' pd='96u*2+14u' ps='96u*2+14u'
m5 z b n1 vss n w=93u l=2.3636u ad='93u*5u+12p' as='93u*5u+12p' pd='93u*2+14u' ps='93u*2+14u'
m6 z a2 n2 vdd p w=217u l=2.3636u ad='217u*5u+12p' as='217u*5u+12p' pd='217u*2+14u' ps='217u*2+14u'
.ends
