* Spice description of noa3ao322_x4
* Spice driver version 134999461
* Date 31/05/2007 at 10:39:14
* ssxlib 0.13um values
.subckt noa3ao322_x4 i0 i1 i2 i3 i4 i5 i6 nq vdd vss
Mtr_00001 vss   sig1  nq    vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00002 nq    sig1  vss   vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00003 sig1  sig4  vss   vss n  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
Mtr_00004 vss   i5    sig8  vss n  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
Mtr_00005 vss   i3    sig8  vss n  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
Mtr_00006 sig5  i0    vss   vss n  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
Mtr_00007 sig4  i2    sig9  vss n  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
Mtr_00008 sig8  i4    vss   vss n  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
Mtr_00009 sig9  i1    sig5  vss n  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
Mtr_00010 sig8  i6    sig4  vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
Mtr_00011 vdd   sig4  sig1  vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
Mtr_00012 vdd   i1    sig16 vdd p  L=0.12U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U
Mtr_00013 sig16 i5    sig17 vdd p  L=0.12U  W=1.65U  AS=0.43725P  AD=0.43725P  PS=3.83U   PD=3.83U
Mtr_00014 sig17 i4    sig18 vdd p  L=0.12U  W=1.595U AS=0.422675P AD=0.422675P PS=3.72U   PD=3.72U
Mtr_00015 sig16 i0    vdd   vdd p  L=0.12U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U
Mtr_00016 nq    sig1  vdd   vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
Mtr_00017 sig16 i2    vdd   vdd p  L=0.12U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U
Mtr_00018 sig4  i6    sig16 vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
Mtr_00019 vdd   sig1  nq    vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
Mtr_00020 sig18 i3    sig4  vdd p  L=0.12U  W=1.595U AS=0.422675P AD=0.422675P PS=3.72U   PD=3.72U
C6  i0    vss   0.654f
C7  i1    vss   0.639f
C10 i2    vss   0.532f
C13 i3    vss   0.654f
C14 i4    vss   0.647f
C12 i5    vss   0.639f
C11 i6    vss   0.575f
C3  nq    vss   0.771f
C1  sig1  vss   0.792f
C16 sig16 vss   0.463f
C4  sig4  vss   1.058f
C8  sig8  vss   0.198f
.ends
