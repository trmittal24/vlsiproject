* Spice description of oai21_x1
* Spice driver version 134934782
* Date 15/09/2003 at 17:05:10
*
.subckt oai21_x1 a1 a2 b vdd vss z 
M3  vdd   b     z     vdd p  L=0.13U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U  
M1  sig5  a1    vdd   vdd p  L=0.13U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U  
M2  z     a2    sig5  vdd p  L=0.13U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U  
M6  sig1  b     z     vss n  L=0.13U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U  
M4  sig1  a1    vss   vss n  L=0.13U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U  
M5  vss   a2    sig1  vss n  L=0.13U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U  
C8  a2    vss   1.549f
C7  b     vss   1.638f
C6  a1    vss   0.989f
C4  vdd   vss   1.059f
C2  z     vss   2.536f
C1  sig1  vss   0.529f
.ends
